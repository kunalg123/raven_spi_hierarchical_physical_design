magic
tech scmos
timestamp 1560666112
<< metal1 >>
rect 960 1303 962 1307
rect 966 1303 969 1307
rect 973 1303 976 1307
rect 966 1288 974 1291
rect 734 1272 737 1281
rect 42 1268 49 1271
rect 706 1268 713 1271
rect 446 1238 470 1241
rect 1422 1238 1430 1241
rect 440 1203 442 1207
rect 446 1203 449 1207
rect 453 1203 456 1207
rect 293 1188 294 1192
rect 354 1188 355 1192
rect 629 1188 630 1192
rect 874 1188 875 1192
rect 717 1168 718 1172
rect 278 1151 281 1161
rect 262 1148 281 1151
rect 294 1148 321 1151
rect 326 1148 334 1151
rect 366 1151 369 1161
rect 366 1148 385 1151
rect 575 1148 582 1151
rect 614 1151 617 1161
rect 598 1148 617 1151
rect 630 1148 657 1151
rect 702 1151 705 1161
rect 762 1158 769 1161
rect 778 1158 782 1162
rect 666 1148 681 1151
rect 686 1148 705 1151
rect 718 1148 726 1151
rect 738 1148 745 1151
rect 750 1148 766 1151
rect 782 1148 790 1151
rect 822 1151 825 1161
rect 822 1148 841 1151
rect 886 1148 918 1151
rect 1102 1148 1113 1151
rect 390 1138 398 1141
rect 678 1138 681 1148
rect 846 1138 849 1148
rect 1126 1138 1134 1141
rect 1134 1128 1153 1131
rect 1162 1128 1177 1131
rect 1430 1118 1438 1121
rect 960 1103 962 1107
rect 966 1103 969 1107
rect 973 1103 976 1107
rect 730 1078 737 1081
rect 183 1068 201 1071
rect 306 1068 313 1071
rect 342 1062 345 1071
rect 390 1068 398 1071
rect 614 1068 622 1071
rect 654 1068 665 1071
rect 1038 1071 1041 1081
rect 1038 1068 1057 1071
rect 206 1058 225 1061
rect 262 1058 278 1061
rect 314 1058 321 1061
rect 350 1058 369 1061
rect 410 1058 425 1061
rect 1126 1058 1145 1061
rect 1327 1058 1345 1061
rect 182 1048 190 1051
rect 222 1048 225 1058
rect 278 1048 281 1058
rect 366 1048 369 1058
rect 686 1048 697 1051
rect 1126 1052 1129 1058
rect 958 1048 966 1051
rect 1430 1038 1441 1041
rect 1438 1032 1441 1038
rect 440 1003 442 1007
rect 446 1003 449 1007
rect 453 1003 456 1007
rect 370 988 371 992
rect 394 988 395 992
rect 794 988 795 992
rect 986 988 993 991
rect 166 948 169 958
rect 398 948 406 951
rect 422 948 441 951
rect 918 948 937 951
rect 422 942 425 948
rect 502 938 510 941
rect 778 938 785 941
rect 902 938 910 941
rect 354 928 361 931
rect 466 928 473 931
rect 510 928 529 931
rect 949 928 950 932
rect 960 903 962 907
rect 966 903 969 907
rect 973 903 976 907
rect 1138 888 1145 891
rect 198 878 214 881
rect 230 872 233 881
rect 374 878 398 881
rect 882 878 889 881
rect 22 868 30 871
rect 250 868 257 871
rect 758 868 774 871
rect 790 868 809 871
rect 894 868 905 871
rect 1158 868 1166 871
rect 238 858 257 861
rect 294 858 302 861
rect 334 861 337 868
rect 326 858 337 861
rect 858 858 886 861
rect 894 858 905 861
rect 934 858 966 861
rect 998 858 1006 861
rect 1062 858 1078 861
rect 1418 858 1425 861
rect 902 852 905 858
rect 1070 848 1078 851
rect 1226 848 1230 852
rect 366 838 390 841
rect 440 803 442 807
rect 446 803 449 807
rect 453 803 456 807
rect 101 788 102 792
rect 741 788 742 792
rect 442 778 443 782
rect 958 768 1001 771
rect 926 766 930 768
rect 126 758 134 761
rect 926 758 937 761
rect 1154 758 1161 761
rect 838 752 842 754
rect 198 748 217 751
rect 534 748 553 751
rect 974 751 978 754
rect 974 748 990 751
rect 910 738 913 748
rect 1022 738 1041 741
rect 1022 732 1025 738
rect 229 728 230 732
rect 1014 728 1022 731
rect 1194 728 1201 731
rect 960 703 962 707
rect 966 703 969 707
rect 973 703 976 707
rect 178 678 185 681
rect 846 678 857 681
rect 218 668 225 671
rect 846 668 857 671
rect 1002 668 1009 671
rect 1038 668 1046 671
rect 1082 668 1089 671
rect 1094 668 1129 671
rect 206 658 225 661
rect 438 658 481 661
rect 518 661 521 668
rect 854 662 857 668
rect 518 658 545 661
rect 610 658 617 661
rect 958 658 985 661
rect 1054 658 1062 661
rect 982 648 1001 651
rect 1018 648 1025 651
rect 630 638 638 641
rect 1430 638 1438 641
rect 618 618 619 622
rect 440 603 442 607
rect 446 603 449 607
rect 453 603 456 607
rect 658 568 665 571
rect 1110 568 1121 571
rect 1110 562 1113 568
rect 1158 561 1162 564
rect 1154 558 1162 561
rect 186 548 193 551
rect 718 548 726 551
rect 1046 548 1065 551
rect 1142 551 1146 554
rect 1138 548 1146 551
rect 186 538 193 541
rect 402 538 409 541
rect 702 538 705 548
rect 726 538 745 541
rect 1018 538 1041 541
rect 1150 531 1153 538
rect 1150 528 1161 531
rect 1182 528 1190 531
rect 426 518 428 522
rect 960 503 962 507
rect 966 503 969 507
rect 973 503 976 507
rect 962 488 963 492
rect 610 478 612 482
rect 854 478 865 481
rect 1338 478 1345 481
rect 414 468 425 471
rect 558 468 585 471
rect 1122 468 1134 471
rect 1142 468 1150 471
rect 1158 468 1166 471
rect 1178 468 1185 471
rect 1198 468 1209 471
rect 1298 468 1313 471
rect 158 458 161 468
rect 422 462 425 468
rect 1198 462 1201 468
rect 510 458 526 461
rect 542 458 550 461
rect 686 458 713 461
rect 910 458 918 461
rect 986 458 993 461
rect 1010 458 1018 461
rect 1222 461 1225 468
rect 1222 458 1233 461
rect 1310 458 1313 468
rect 1318 458 1337 461
rect 1014 456 1018 458
rect 614 438 630 441
rect 1430 438 1438 441
rect 538 418 539 422
rect 714 418 715 422
rect 440 403 442 407
rect 446 403 449 407
rect 453 403 456 407
rect 602 388 603 392
rect 1014 372 1017 381
rect 199 348 206 351
rect 518 348 537 351
rect 854 348 865 351
rect 862 342 865 348
rect 1086 351 1090 352
rect 1166 351 1169 361
rect 1074 348 1090 351
rect 1150 348 1169 351
rect 1194 348 1201 351
rect 402 338 409 341
rect 454 338 486 341
rect 682 338 689 341
rect 878 341 881 348
rect 870 338 881 341
rect 1070 338 1073 348
rect 1102 338 1110 341
rect 1190 338 1193 348
rect 1422 338 1438 341
rect 418 328 430 331
rect 626 328 630 332
rect 774 321 777 328
rect 766 318 777 321
rect 960 303 962 307
rect 966 303 969 307
rect 973 303 976 307
rect 794 288 795 292
rect 343 268 361 271
rect 430 268 438 271
rect 502 271 505 281
rect 518 278 537 281
rect 614 278 622 281
rect 1002 278 1014 281
rect 446 268 489 271
rect 502 268 521 271
rect 978 268 993 271
rect 1010 268 1025 271
rect 126 258 129 268
rect 374 261 377 268
rect 366 258 377 261
rect 622 258 630 261
rect 822 251 825 258
rect 822 248 833 251
rect 918 248 945 251
rect 538 238 545 241
rect 966 218 982 221
rect 440 203 442 207
rect 446 203 449 207
rect 453 203 456 207
rect 634 188 635 192
rect 1186 188 1187 192
rect 574 158 593 161
rect 962 158 966 162
rect 986 158 1001 161
rect 1066 158 1070 162
rect 1218 158 1222 162
rect 286 148 329 151
rect 390 148 398 151
rect 458 148 473 151
rect 606 148 614 151
rect 294 138 310 141
rect 338 138 345 141
rect 414 138 422 141
rect 442 138 462 141
rect 534 141 537 148
rect 638 142 641 151
rect 734 148 742 151
rect 798 151 802 152
rect 798 148 806 151
rect 810 148 814 151
rect 974 148 1009 151
rect 1022 148 1033 151
rect 1082 148 1089 151
rect 1166 148 1177 151
rect 526 138 537 141
rect 694 138 702 141
rect 922 138 929 141
rect 974 138 977 148
rect 1022 138 1025 148
rect 1030 142 1033 148
rect 1094 138 1110 141
rect 1174 138 1177 148
rect 822 128 841 131
rect 1046 128 1049 138
rect 1246 128 1254 131
rect 517 118 518 122
rect 960 103 962 107
rect 966 103 969 107
rect 973 103 976 107
rect 394 88 401 91
rect 933 88 934 92
rect 262 78 278 81
rect 286 78 305 81
rect 338 78 345 81
rect 438 78 446 81
rect 590 78 598 82
rect 714 78 726 81
rect 1146 78 1161 81
rect 590 72 593 78
rect 306 68 313 71
rect 610 68 625 71
rect 974 68 982 71
rect 1054 68 1065 71
rect 1126 71 1129 78
rect 1126 68 1137 71
rect 518 58 534 61
rect 554 58 561 61
rect 662 58 670 61
rect 910 58 929 61
rect 1098 58 1105 61
rect 1338 58 1345 61
rect 1382 58 1390 61
rect 382 48 390 51
rect 586 48 593 51
rect 926 48 929 58
rect 974 51 977 58
rect 974 48 1001 51
rect 440 3 442 7
rect 446 3 449 7
rect 453 3 456 7
<< m2contact >>
rect 962 1303 966 1307
rect 969 1303 973 1307
rect 262 1288 266 1292
rect 494 1288 498 1292
rect 926 1288 930 1292
rect 974 1288 978 1292
rect 1182 1288 1186 1292
rect 1206 1288 1210 1292
rect 1254 1288 1258 1292
rect 1278 1288 1282 1292
rect 1302 1288 1306 1292
rect 1326 1288 1330 1292
rect 1374 1288 1378 1292
rect 174 1278 178 1282
rect 366 1278 370 1282
rect 614 1278 618 1282
rect 758 1278 762 1282
rect 838 1278 842 1282
rect 1078 1278 1082 1282
rect 1174 1279 1178 1283
rect 1198 1279 1202 1283
rect 1222 1279 1226 1283
rect 1230 1278 1234 1282
rect 1246 1279 1250 1283
rect 1270 1279 1274 1283
rect 1294 1279 1298 1283
rect 1366 1279 1370 1283
rect 1390 1279 1394 1283
rect 1414 1279 1418 1283
rect 6 1268 10 1272
rect 38 1268 42 1272
rect 190 1268 194 1272
rect 350 1268 354 1272
rect 502 1268 506 1272
rect 630 1268 634 1272
rect 702 1268 706 1272
rect 734 1268 738 1272
rect 854 1268 858 1272
rect 1094 1268 1098 1272
rect 62 1258 66 1262
rect 230 1258 234 1262
rect 278 1258 282 1262
rect 302 1258 306 1262
rect 406 1258 410 1262
rect 478 1258 482 1262
rect 518 1258 522 1262
rect 574 1258 578 1262
rect 678 1258 682 1262
rect 726 1258 730 1262
rect 798 1258 802 1262
rect 942 1258 946 1262
rect 950 1258 954 1262
rect 1038 1258 1042 1262
rect 1134 1258 1138 1262
rect 1166 1258 1170 1262
rect 1190 1258 1194 1262
rect 1214 1258 1218 1262
rect 1238 1258 1242 1262
rect 1262 1258 1266 1262
rect 1286 1258 1290 1262
rect 1310 1258 1314 1262
rect 1334 1258 1338 1262
rect 1358 1258 1362 1262
rect 1382 1258 1386 1262
rect 1406 1258 1410 1262
rect 238 1248 242 1252
rect 302 1248 306 1252
rect 678 1248 682 1252
rect 902 1248 906 1252
rect 1142 1248 1146 1252
rect 470 1238 474 1242
rect 1318 1238 1322 1242
rect 1430 1238 1434 1242
rect 798 1227 802 1231
rect 14 1218 18 1222
rect 94 1218 98 1222
rect 238 1218 242 1222
rect 302 1218 306 1222
rect 534 1218 538 1222
rect 678 1218 682 1222
rect 742 1218 746 1222
rect 998 1218 1002 1222
rect 1142 1218 1146 1222
rect 1350 1218 1354 1222
rect 1398 1218 1402 1222
rect 1366 1208 1370 1212
rect 1390 1208 1394 1212
rect 1414 1208 1418 1212
rect 442 1203 446 1207
rect 449 1203 453 1207
rect 1334 1198 1338 1202
rect 30 1188 34 1192
rect 70 1188 74 1192
rect 294 1188 298 1192
rect 350 1188 354 1192
rect 630 1188 634 1192
rect 870 1188 874 1192
rect 1358 1188 1362 1192
rect 182 1178 186 1182
rect 446 1179 450 1183
rect 1054 1179 1058 1183
rect 1270 1178 1274 1182
rect 718 1168 722 1172
rect 214 1156 218 1160
rect 230 1158 234 1162
rect 270 1158 274 1162
rect 22 1148 26 1152
rect 46 1148 50 1152
rect 54 1148 58 1152
rect 85 1148 89 1152
rect 182 1148 186 1152
rect 310 1158 314 1162
rect 334 1148 338 1152
rect 350 1148 354 1152
rect 374 1158 378 1162
rect 446 1156 450 1160
rect 606 1158 610 1162
rect 430 1148 434 1152
rect 582 1148 586 1152
rect 646 1158 650 1162
rect 694 1158 698 1162
rect 662 1148 666 1152
rect 758 1158 762 1162
rect 782 1158 786 1162
rect 726 1148 730 1152
rect 734 1148 738 1152
rect 766 1148 770 1152
rect 790 1148 794 1152
rect 806 1148 810 1152
rect 830 1158 834 1162
rect 1054 1156 1058 1160
rect 1302 1156 1306 1160
rect 846 1148 850 1152
rect 854 1148 858 1152
rect 862 1148 866 1152
rect 918 1148 922 1152
rect 966 1148 970 1152
rect 1142 1148 1146 1152
rect 1270 1148 1274 1152
rect 1342 1148 1346 1152
rect 1366 1148 1370 1152
rect 1390 1148 1394 1152
rect 1414 1148 1418 1152
rect 6 1138 10 1142
rect 182 1138 186 1142
rect 254 1138 258 1142
rect 302 1138 306 1142
rect 334 1138 338 1142
rect 342 1138 346 1142
rect 398 1138 402 1142
rect 478 1138 482 1142
rect 590 1138 594 1142
rect 638 1138 642 1142
rect 670 1138 674 1142
rect 726 1138 730 1142
rect 734 1138 738 1142
rect 790 1138 794 1142
rect 798 1138 802 1142
rect 925 1138 929 1142
rect 1022 1138 1026 1142
rect 1118 1138 1122 1142
rect 1134 1138 1138 1142
rect 1270 1138 1274 1142
rect 1406 1138 1410 1142
rect 166 1128 170 1132
rect 494 1128 498 1132
rect 822 1128 826 1132
rect 1006 1128 1010 1132
rect 1094 1128 1098 1132
rect 1158 1128 1162 1132
rect 1254 1128 1258 1132
rect 1382 1118 1386 1122
rect 1438 1118 1442 1122
rect 962 1103 966 1107
rect 969 1103 973 1107
rect 630 1088 634 1092
rect 758 1088 762 1092
rect 1006 1088 1010 1092
rect 1030 1088 1034 1092
rect 1358 1088 1362 1092
rect 1406 1088 1410 1092
rect 14 1078 18 1082
rect 102 1078 106 1082
rect 222 1078 226 1082
rect 502 1078 506 1082
rect 638 1078 642 1082
rect 646 1078 650 1082
rect 686 1078 690 1082
rect 726 1078 730 1082
rect 742 1078 746 1082
rect 766 1078 770 1082
rect 862 1078 866 1082
rect 86 1068 90 1072
rect 246 1068 250 1072
rect 270 1068 274 1072
rect 278 1068 282 1072
rect 302 1068 306 1072
rect 326 1068 330 1072
rect 374 1068 378 1072
rect 398 1068 402 1072
rect 518 1068 522 1072
rect 590 1068 594 1072
rect 622 1068 626 1072
rect 878 1068 882 1072
rect 966 1068 970 1072
rect 1022 1068 1026 1072
rect 1046 1078 1050 1082
rect 1246 1078 1250 1082
rect 1374 1079 1378 1083
rect 1078 1068 1082 1072
rect 1094 1068 1098 1072
rect 1110 1068 1114 1072
rect 1134 1068 1138 1072
rect 1158 1068 1162 1072
rect 1230 1068 1234 1072
rect 46 1058 50 1062
rect 142 1058 146 1062
rect 238 1058 242 1062
rect 278 1058 282 1062
rect 294 1058 298 1062
rect 310 1058 314 1062
rect 342 1058 346 1062
rect 382 1058 386 1062
rect 406 1058 410 1062
rect 550 1058 554 1062
rect 574 1058 578 1062
rect 606 1058 610 1062
rect 622 1058 626 1062
rect 670 1058 674 1062
rect 710 1058 714 1062
rect 726 1058 730 1062
rect 750 1058 754 1062
rect 822 1058 826 1062
rect 934 1058 938 1062
rect 990 1058 994 1062
rect 1014 1058 1018 1062
rect 1062 1058 1066 1062
rect 1070 1058 1074 1062
rect 1102 1058 1106 1062
rect 1118 1058 1122 1062
rect 1190 1058 1194 1062
rect 1286 1058 1290 1062
rect 1366 1058 1370 1062
rect 1390 1058 1394 1062
rect 1414 1058 1418 1062
rect 38 1048 42 1052
rect 190 1048 194 1052
rect 214 1048 218 1052
rect 334 1048 338 1052
rect 358 1048 362 1052
rect 566 1048 570 1052
rect 590 1048 594 1052
rect 718 1048 722 1052
rect 910 1050 914 1054
rect 950 1048 954 1052
rect 966 1048 970 1052
rect 1126 1048 1130 1052
rect 1158 1048 1162 1052
rect 1198 1050 1202 1054
rect 702 1038 706 1042
rect 782 1038 786 1042
rect 910 1027 914 1031
rect 1198 1027 1202 1031
rect 1438 1028 1442 1032
rect 6 1018 10 1022
rect 38 1018 42 1022
rect 566 1018 570 1022
rect 1094 1018 1098 1022
rect 1326 1018 1330 1022
rect 1382 1018 1386 1022
rect 442 1003 446 1007
rect 449 1003 453 1007
rect 1414 998 1418 1002
rect 14 988 18 992
rect 158 988 162 992
rect 198 988 202 992
rect 366 988 370 992
rect 390 988 394 992
rect 406 988 410 992
rect 438 988 442 992
rect 478 988 482 992
rect 790 988 794 992
rect 830 988 834 992
rect 862 988 866 992
rect 982 988 986 992
rect 1038 988 1042 992
rect 1230 988 1234 992
rect 1406 988 1410 992
rect 1438 988 1442 992
rect 606 978 610 982
rect 1134 978 1138 982
rect 1278 979 1282 983
rect 702 968 706 972
rect 838 968 842 972
rect 870 968 874 972
rect 894 968 898 972
rect 1046 968 1050 972
rect 158 958 162 962
rect 166 958 170 962
rect 198 958 202 962
rect 558 958 562 962
rect 726 958 730 962
rect 822 958 826 962
rect 854 958 858 962
rect 886 958 890 962
rect 1062 958 1066 962
rect 1086 958 1090 962
rect 54 948 58 952
rect 1278 956 1282 960
rect 198 948 202 952
rect 302 948 306 952
rect 374 948 378 952
rect 406 948 410 952
rect 486 948 490 952
rect 518 948 522 952
rect 606 948 610 952
rect 718 948 722 952
rect 750 948 754 952
rect 766 948 770 952
rect 790 948 794 952
rect 806 948 810 952
rect 830 948 834 952
rect 862 948 866 952
rect 958 948 962 952
rect 966 948 970 952
rect 1014 948 1018 952
rect 1030 948 1034 952
rect 1054 948 1058 952
rect 1134 948 1138 952
rect 1262 948 1266 952
rect 1422 948 1426 952
rect 110 938 114 942
rect 246 938 250 942
rect 422 938 426 942
rect 430 938 434 942
rect 494 938 498 942
rect 510 938 514 942
rect 606 938 610 942
rect 742 938 746 942
rect 758 938 762 942
rect 774 938 778 942
rect 814 938 818 942
rect 910 938 914 942
rect 1022 938 1026 942
rect 1134 938 1138 942
rect 1310 938 1314 942
rect 94 928 98 932
rect 262 928 266 932
rect 350 928 354 932
rect 382 928 386 932
rect 422 928 426 932
rect 462 928 466 932
rect 534 928 538 932
rect 622 928 626 932
rect 734 928 738 932
rect 910 928 914 932
rect 950 928 954 932
rect 998 928 1002 932
rect 1006 928 1010 932
rect 1150 928 1154 932
rect 1326 928 1330 932
rect 342 918 346 922
rect 1230 918 1234 922
rect 962 903 966 907
rect 969 903 973 907
rect 318 888 322 892
rect 358 888 362 892
rect 734 888 738 892
rect 782 888 786 892
rect 806 888 810 892
rect 862 888 866 892
rect 918 888 922 892
rect 1006 888 1010 892
rect 1118 888 1122 892
rect 1134 888 1138 892
rect 1414 888 1418 892
rect 1438 888 1442 892
rect 118 878 122 882
rect 214 878 218 882
rect 302 878 306 882
rect 310 878 314 882
rect 398 878 402 882
rect 486 878 490 882
rect 654 878 658 882
rect 798 878 802 882
rect 870 878 874 882
rect 878 878 882 882
rect 942 878 946 882
rect 1014 878 1018 882
rect 1038 878 1042 882
rect 1126 878 1130 882
rect 1166 878 1170 882
rect 1326 878 1330 882
rect 30 868 34 872
rect 102 868 106 872
rect 230 868 234 872
rect 246 868 250 872
rect 334 868 338 872
rect 502 868 506 872
rect 638 868 642 872
rect 750 868 754 872
rect 774 868 778 872
rect 862 868 866 872
rect 1006 868 1010 872
rect 1030 868 1034 872
rect 1054 868 1058 872
rect 1118 868 1122 872
rect 1166 868 1170 872
rect 1174 868 1178 872
rect 1190 868 1194 872
rect 1206 868 1210 872
rect 1238 868 1242 872
rect 1310 868 1314 872
rect 6 858 10 862
rect 54 858 58 862
rect 278 858 282 862
rect 286 858 290 862
rect 302 858 306 862
rect 342 858 346 862
rect 550 858 554 862
rect 590 858 594 862
rect 814 858 818 862
rect 854 858 858 862
rect 886 858 890 862
rect 926 858 930 862
rect 966 858 970 862
rect 1006 858 1010 862
rect 1078 858 1082 862
rect 1110 858 1114 862
rect 1198 858 1202 862
rect 1230 858 1234 862
rect 1262 858 1266 862
rect 1407 858 1411 862
rect 1414 858 1418 862
rect 54 848 58 852
rect 358 848 362 852
rect 534 850 538 854
rect 606 850 610 854
rect 766 848 770 852
rect 902 848 906 852
rect 918 848 922 852
rect 1046 848 1050 852
rect 1078 848 1082 852
rect 1142 848 1146 852
rect 1182 848 1186 852
rect 1214 848 1218 852
rect 1230 848 1234 852
rect 1278 850 1282 854
rect 390 838 394 842
rect 534 827 538 831
rect 606 827 610 831
rect 1278 827 1282 831
rect 54 818 58 822
rect 222 818 226 822
rect 406 818 410 822
rect 442 803 446 807
rect 449 803 453 807
rect 62 788 66 792
rect 102 788 106 792
rect 158 788 162 792
rect 414 788 418 792
rect 478 788 482 792
rect 558 788 562 792
rect 646 788 650 792
rect 678 788 682 792
rect 742 788 746 792
rect 774 788 778 792
rect 830 788 834 792
rect 862 788 866 792
rect 886 788 890 792
rect 966 788 970 792
rect 1070 788 1074 792
rect 1110 788 1114 792
rect 1142 788 1146 792
rect 1182 788 1186 792
rect 1238 788 1242 792
rect 286 779 290 783
rect 438 778 442 782
rect 1390 779 1394 783
rect 766 768 770 772
rect 822 768 826 772
rect 854 768 858 772
rect 894 768 898 772
rect 926 768 930 772
rect 1134 768 1138 772
rect 1174 768 1178 772
rect 134 758 138 762
rect 286 756 290 760
rect 454 758 458 762
rect 710 758 714 762
rect 726 758 730 762
rect 782 758 786 762
rect 870 758 874 762
rect 878 758 882 762
rect 1102 758 1106 762
rect 1150 758 1154 762
rect 1390 756 1394 760
rect 86 748 90 752
rect 110 748 114 752
rect 118 748 122 752
rect 150 748 154 752
rect 174 748 178 752
rect 182 748 186 752
rect 238 748 242 752
rect 246 748 250 752
rect 270 748 274 752
rect 438 748 442 752
rect 518 748 522 752
rect 574 748 578 752
rect 582 748 586 752
rect 670 748 674 752
rect 694 748 698 752
rect 702 748 706 752
rect 742 748 746 752
rect 774 748 778 752
rect 790 748 794 752
rect 830 748 834 752
rect 838 748 842 752
rect 862 748 866 752
rect 886 748 890 752
rect 910 748 914 752
rect 966 748 970 752
rect 990 748 994 752
rect 998 748 1002 752
rect 1046 748 1050 752
rect 1094 748 1098 752
rect 1142 748 1146 752
rect 1166 748 1170 752
rect 1214 748 1218 752
rect 1398 748 1402 752
rect 6 738 10 742
rect 318 738 322 742
rect 430 738 434 742
rect 590 738 594 742
rect 750 738 754 742
rect 798 738 802 742
rect 1086 738 1090 742
rect 1118 738 1122 742
rect 1206 738 1210 742
rect 1358 738 1362 742
rect 134 728 138 732
rect 190 728 194 732
rect 230 728 234 732
rect 334 728 338 732
rect 486 728 490 732
rect 526 728 530 732
rect 718 728 722 732
rect 806 728 810 732
rect 942 728 946 732
rect 1022 728 1026 732
rect 1030 728 1034 732
rect 1190 728 1194 732
rect 1342 728 1346 732
rect 502 718 506 722
rect 534 718 538 722
rect 926 718 930 722
rect 1262 718 1266 722
rect 962 703 966 707
rect 969 703 973 707
rect 166 688 170 692
rect 422 688 426 692
rect 814 688 818 692
rect 886 688 890 692
rect 910 688 914 692
rect 950 688 954 692
rect 1022 688 1026 692
rect 1070 688 1074 692
rect 1126 688 1130 692
rect 1190 688 1194 692
rect 86 678 90 682
rect 174 678 178 682
rect 190 678 194 682
rect 198 678 202 682
rect 342 678 346 682
rect 446 678 450 682
rect 518 678 522 682
rect 726 678 730 682
rect 838 678 842 682
rect 894 678 898 682
rect 902 678 906 682
rect 942 678 946 682
rect 990 678 994 682
rect 1046 678 1050 682
rect 1078 678 1082 682
rect 1118 678 1122 682
rect 1182 678 1186 682
rect 1326 678 1330 682
rect 70 668 74 672
rect 214 668 218 672
rect 326 668 330 672
rect 518 668 522 672
rect 598 668 602 672
rect 606 668 610 672
rect 742 668 746 672
rect 830 668 834 672
rect 926 668 930 672
rect 998 668 1002 672
rect 1014 668 1018 672
rect 1046 668 1050 672
rect 1078 668 1082 672
rect 1190 668 1194 672
rect 1342 668 1346 672
rect 38 658 42 662
rect 246 658 250 662
rect 254 658 258 662
rect 294 658 298 662
rect 502 658 506 662
rect 510 658 514 662
rect 566 658 570 662
rect 574 658 578 662
rect 606 658 610 662
rect 686 658 690 662
rect 782 658 786 662
rect 854 658 858 662
rect 870 658 874 662
rect 878 658 882 662
rect 918 658 922 662
rect 1062 658 1066 662
rect 1134 658 1138 662
rect 1198 658 1202 662
rect 1286 658 1290 662
rect 1398 658 1402 662
rect 1414 658 1418 662
rect 22 648 26 652
rect 278 648 282 652
rect 550 648 554 652
rect 774 650 778 654
rect 814 648 818 652
rect 862 648 866 652
rect 1014 648 1018 652
rect 1102 648 1106 652
rect 1374 650 1378 654
rect 638 638 642 642
rect 934 638 938 642
rect 1438 638 1442 642
rect 774 627 778 631
rect 1374 627 1378 631
rect 22 618 26 622
rect 182 618 186 622
rect 278 618 282 622
rect 438 618 442 622
rect 486 618 490 622
rect 590 618 594 622
rect 614 618 618 622
rect 646 618 650 622
rect 1246 618 1250 622
rect 442 603 446 607
rect 449 603 453 607
rect 22 588 26 592
rect 166 588 170 592
rect 246 588 250 592
rect 390 588 394 592
rect 494 588 498 592
rect 638 588 642 592
rect 854 588 858 592
rect 998 588 1002 592
rect 1174 588 1178 592
rect 1342 588 1346 592
rect 654 568 658 572
rect 22 558 26 562
rect 246 558 250 562
rect 494 558 498 562
rect 694 558 698 562
rect 702 558 706 562
rect 734 558 738 562
rect 774 558 778 562
rect 806 558 810 562
rect 830 558 834 562
rect 854 558 858 562
rect 1054 558 1058 562
rect 1110 558 1114 562
rect 1150 558 1154 562
rect 1342 558 1346 562
rect 22 548 26 552
rect 38 548 42 552
rect 182 548 186 552
rect 214 548 218 552
rect 222 548 226 552
rect 246 548 250 552
rect 294 548 298 552
rect 502 548 506 552
rect 678 548 682 552
rect 686 548 690 552
rect 702 548 706 552
rect 726 548 730 552
rect 790 548 794 552
rect 798 548 802 552
rect 862 548 866 552
rect 1070 548 1074 552
rect 1102 548 1106 552
rect 1118 548 1122 552
rect 1134 548 1138 552
rect 1158 548 1162 552
rect 1294 548 1298 552
rect 70 538 74 542
rect 182 538 186 542
rect 294 538 298 542
rect 398 538 402 542
rect 542 538 546 542
rect 670 538 674 542
rect 750 538 754 542
rect 758 538 762 542
rect 782 538 786 542
rect 814 538 818 542
rect 902 538 906 542
rect 1014 538 1018 542
rect 1078 538 1082 542
rect 1110 538 1114 542
rect 1150 538 1154 542
rect 1197 538 1201 542
rect 1294 538 1298 542
rect 1366 538 1370 542
rect 1430 538 1434 542
rect 86 528 90 532
rect 310 528 314 532
rect 558 528 562 532
rect 654 528 658 532
rect 918 528 922 532
rect 1030 528 1034 532
rect 1134 528 1138 532
rect 1190 528 1194 532
rect 1278 528 1282 532
rect 422 518 426 522
rect 774 518 778 522
rect 830 518 834 522
rect 1086 518 1090 522
rect 962 503 966 507
rect 969 503 973 507
rect 22 488 26 492
rect 438 488 442 492
rect 590 488 594 492
rect 662 488 666 492
rect 750 488 754 492
rect 782 488 786 492
rect 798 488 802 492
rect 806 488 810 492
rect 870 488 874 492
rect 958 488 962 492
rect 1222 488 1226 492
rect 1254 488 1258 492
rect 1286 488 1290 492
rect 1382 488 1386 492
rect 118 478 122 482
rect 294 478 298 482
rect 446 478 450 482
rect 526 478 530 482
rect 550 478 554 482
rect 598 478 602 482
rect 606 478 610 482
rect 654 478 658 482
rect 942 478 946 482
rect 1006 478 1010 482
rect 1046 478 1050 482
rect 1102 478 1106 482
rect 1134 478 1138 482
rect 1174 478 1178 482
rect 1246 478 1250 482
rect 1278 478 1282 482
rect 1326 478 1330 482
rect 1334 478 1338 482
rect 1350 478 1354 482
rect 102 468 106 472
rect 158 468 162 472
rect 278 468 282 472
rect 398 468 402 472
rect 430 468 434 472
rect 470 468 474 472
rect 486 468 490 472
rect 502 468 506 472
rect 518 468 522 472
rect 638 468 642 472
rect 646 468 650 472
rect 678 468 682 472
rect 702 468 706 472
rect 734 468 738 472
rect 758 468 762 472
rect 790 468 794 472
rect 822 468 826 472
rect 830 468 834 472
rect 878 468 882 472
rect 902 468 906 472
rect 918 468 922 472
rect 934 468 938 472
rect 950 468 954 472
rect 1118 468 1122 472
rect 1134 468 1138 472
rect 1150 468 1154 472
rect 1166 468 1170 472
rect 1174 468 1178 472
rect 1190 468 1194 472
rect 1222 468 1226 472
rect 1238 468 1242 472
rect 1262 468 1266 472
rect 1294 468 1298 472
rect 1358 468 1362 472
rect 1406 468 1410 472
rect 6 458 10 462
rect 54 458 58 462
rect 230 458 234 462
rect 406 458 410 462
rect 422 458 426 462
rect 478 458 482 462
rect 494 458 498 462
rect 526 458 530 462
rect 550 458 554 462
rect 566 458 570 462
rect 574 458 578 462
rect 622 458 626 462
rect 670 458 674 462
rect 766 458 770 462
rect 838 458 842 462
rect 886 458 890 462
rect 918 458 922 462
rect 926 458 930 462
rect 982 458 986 462
rect 1006 458 1010 462
rect 1022 458 1026 462
rect 1062 458 1066 462
rect 1086 458 1090 462
rect 1126 458 1130 462
rect 1198 458 1202 462
rect 1270 458 1274 462
rect 1302 458 1306 462
rect 1414 458 1418 462
rect 54 448 58 452
rect 246 450 250 454
rect 374 448 378 452
rect 390 448 394 452
rect 630 448 634 452
rect 694 448 698 452
rect 726 448 730 452
rect 750 448 754 452
rect 806 448 810 452
rect 854 448 858 452
rect 894 448 898 452
rect 966 448 970 452
rect 998 448 1002 452
rect 1094 448 1098 452
rect 1166 448 1170 452
rect 1222 448 1226 452
rect 1230 448 1234 452
rect 630 438 634 442
rect 1030 438 1034 442
rect 1062 438 1066 442
rect 1078 438 1082 442
rect 1438 438 1442 442
rect 198 428 202 432
rect 246 427 250 431
rect 54 418 58 422
rect 534 418 538 422
rect 710 418 714 422
rect 1038 418 1042 422
rect 1086 418 1090 422
rect 1102 418 1106 422
rect 442 403 446 407
rect 449 403 453 407
rect 54 388 58 392
rect 374 388 378 392
rect 598 388 602 392
rect 926 388 930 392
rect 1126 388 1130 392
rect 1382 388 1386 392
rect 246 379 250 383
rect 574 378 578 382
rect 566 368 570 372
rect 766 368 770 372
rect 798 368 802 372
rect 1014 368 1018 372
rect 1022 368 1026 372
rect 1238 368 1242 372
rect 54 358 58 362
rect 246 356 250 360
rect 422 358 426 362
rect 550 358 554 362
rect 582 358 586 362
rect 654 358 658 362
rect 782 358 786 362
rect 878 358 882 362
rect 910 358 914 362
rect 918 358 922 362
rect 1006 358 1010 362
rect 1158 358 1162 362
rect 6 348 10 352
rect 54 348 58 352
rect 206 348 210 352
rect 230 348 234 352
rect 478 348 482 352
rect 574 348 578 352
rect 606 348 610 352
rect 614 348 618 352
rect 646 348 650 352
rect 702 348 706 352
rect 734 348 738 352
rect 750 348 754 352
rect 774 348 778 352
rect 790 348 794 352
rect 822 348 826 352
rect 878 348 882 352
rect 894 348 898 352
rect 902 348 906 352
rect 974 348 978 352
rect 1014 348 1018 352
rect 1046 348 1050 352
rect 1062 348 1066 352
rect 1070 348 1074 352
rect 1382 358 1386 362
rect 1182 348 1186 352
rect 1190 348 1194 352
rect 1278 348 1282 352
rect 1406 348 1410 352
rect 102 338 106 342
rect 278 338 282 342
rect 398 338 402 342
rect 438 338 442 342
rect 486 338 490 342
rect 526 338 530 342
rect 550 338 554 342
rect 622 338 626 342
rect 638 338 642 342
rect 670 338 674 342
rect 678 338 682 342
rect 694 338 698 342
rect 742 338 746 342
rect 798 338 802 342
rect 814 338 818 342
rect 846 338 850 342
rect 862 338 866 342
rect 886 338 890 342
rect 934 338 938 342
rect 950 338 954 342
rect 1038 338 1042 342
rect 1078 338 1082 342
rect 1110 338 1114 342
rect 1118 338 1122 342
rect 1142 338 1146 342
rect 1174 338 1178 342
rect 1206 338 1210 342
rect 1334 338 1338 342
rect 1438 338 1442 342
rect 118 328 122 332
rect 294 328 298 332
rect 430 328 434 332
rect 502 328 506 332
rect 510 328 514 332
rect 590 328 594 332
rect 622 328 626 332
rect 678 328 682 332
rect 710 328 714 332
rect 726 328 730 332
rect 774 328 778 332
rect 830 328 834 332
rect 1126 328 1130 332
rect 1222 328 1226 332
rect 1318 328 1322 332
rect 22 318 26 322
rect 390 318 394 322
rect 494 318 498 322
rect 654 318 658 322
rect 718 318 722 322
rect 838 318 842 322
rect 942 318 946 322
rect 990 318 994 322
rect 1046 318 1050 322
rect 1214 318 1218 322
rect 962 303 966 307
rect 969 303 973 307
rect 494 288 498 292
rect 678 288 682 292
rect 742 288 746 292
rect 766 288 770 292
rect 790 288 794 292
rect 822 288 826 292
rect 1374 288 1378 292
rect 86 278 90 282
rect 262 278 266 282
rect 390 278 394 282
rect 454 278 458 282
rect 70 268 74 272
rect 126 268 130 272
rect 246 268 250 272
rect 374 268 378 272
rect 398 268 402 272
rect 414 268 418 272
rect 438 268 442 272
rect 510 278 514 282
rect 598 278 602 282
rect 606 278 610 282
rect 622 278 626 282
rect 830 278 834 282
rect 926 278 930 282
rect 1014 278 1018 282
rect 1102 278 1106 282
rect 1278 278 1282 282
rect 550 268 554 272
rect 574 268 578 272
rect 630 268 634 272
rect 694 268 698 272
rect 710 268 714 272
rect 726 268 730 272
rect 782 268 786 272
rect 806 268 810 272
rect 846 268 850 272
rect 870 268 874 272
rect 886 268 890 272
rect 974 268 978 272
rect 1006 268 1010 272
rect 1118 268 1122 272
rect 1294 268 1298 272
rect 1430 268 1434 272
rect 22 258 26 262
rect 198 258 202 262
rect 406 258 410 262
rect 422 258 426 262
rect 438 258 442 262
rect 478 258 482 262
rect 526 258 530 262
rect 558 258 562 262
rect 582 258 586 262
rect 630 258 634 262
rect 638 258 642 262
rect 646 258 650 262
rect 662 258 666 262
rect 702 258 706 262
rect 750 258 754 262
rect 822 258 826 262
rect 854 258 858 262
rect 878 258 882 262
rect 910 258 914 262
rect 950 258 954 262
rect 1062 258 1066 262
rect 1174 258 1178 262
rect 1238 258 1242 262
rect 22 248 26 252
rect 198 248 202 252
rect 574 248 578 252
rect 590 248 594 252
rect 654 248 658 252
rect 718 248 722 252
rect 742 248 746 252
rect 798 248 802 252
rect 862 248 866 252
rect 1006 248 1010 252
rect 1150 250 1154 254
rect 1342 248 1346 252
rect 166 238 170 242
rect 534 238 538 242
rect 902 238 906 242
rect 958 238 962 242
rect 342 228 346 232
rect 1150 227 1154 231
rect 22 218 26 222
rect 198 218 202 222
rect 374 218 378 222
rect 910 218 914 222
rect 982 218 986 222
rect 1198 218 1202 222
rect 1342 218 1346 222
rect 1374 218 1378 222
rect 442 203 446 207
rect 449 203 453 207
rect 62 188 66 192
rect 94 188 98 192
rect 630 188 634 192
rect 662 188 666 192
rect 726 188 730 192
rect 758 188 762 192
rect 854 188 858 192
rect 878 188 882 192
rect 1030 188 1034 192
rect 1182 188 1186 192
rect 1238 188 1242 192
rect 1390 179 1394 183
rect 238 168 242 172
rect 366 168 370 172
rect 94 158 98 162
rect 334 158 338 162
rect 398 158 402 162
rect 478 158 482 162
rect 510 158 514 162
rect 566 158 570 162
rect 950 158 954 162
rect 966 158 970 162
rect 982 158 986 162
rect 1054 158 1058 162
rect 1070 158 1074 162
rect 1134 158 1138 162
rect 1198 158 1202 162
rect 1214 158 1218 162
rect 1230 158 1234 162
rect 1390 156 1394 160
rect 198 148 202 152
rect 350 148 354 152
rect 382 148 386 152
rect 398 148 402 152
rect 446 148 450 152
rect 454 148 458 152
rect 502 148 506 152
rect 534 148 538 152
rect 598 148 602 152
rect 614 148 618 152
rect 6 138 10 142
rect 142 138 146 142
rect 310 138 314 142
rect 318 138 322 142
rect 334 138 338 142
rect 374 138 378 142
rect 422 138 426 142
rect 438 138 442 142
rect 462 138 466 142
rect 478 138 482 142
rect 494 138 498 142
rect 646 148 650 152
rect 678 148 682 152
rect 710 148 714 152
rect 742 148 746 152
rect 806 148 810 152
rect 814 148 818 152
rect 830 148 834 152
rect 854 148 858 152
rect 878 148 882 152
rect 894 148 898 152
rect 910 148 914 152
rect 942 148 946 152
rect 966 148 970 152
rect 1014 148 1018 152
rect 1070 148 1074 152
rect 1078 148 1082 152
rect 1118 148 1122 152
rect 1126 148 1130 152
rect 1150 148 1154 152
rect 1182 148 1186 152
rect 1214 148 1218 152
rect 1261 148 1265 152
rect 1302 148 1306 152
rect 542 138 546 142
rect 582 138 586 142
rect 614 138 618 142
rect 638 138 642 142
rect 702 138 706 142
rect 806 138 810 142
rect 902 138 906 142
rect 918 138 922 142
rect 934 138 938 142
rect 1030 138 1034 142
rect 1046 138 1050 142
rect 1078 138 1082 142
rect 1110 138 1114 142
rect 1142 138 1146 142
rect 1206 138 1210 142
rect 1358 138 1362 142
rect 158 128 162 132
rect 302 128 306 132
rect 406 128 410 132
rect 422 128 426 132
rect 550 128 554 132
rect 558 128 562 132
rect 622 128 626 132
rect 814 128 818 132
rect 862 128 866 132
rect 886 128 890 132
rect 918 128 922 132
rect 1102 128 1106 132
rect 1254 128 1258 132
rect 1342 128 1346 132
rect 294 118 298 122
rect 334 118 338 122
rect 430 118 434 122
rect 518 118 522 122
rect 962 103 966 107
rect 969 103 973 107
rect 86 88 90 92
rect 390 88 394 92
rect 478 88 482 92
rect 502 88 506 92
rect 550 88 554 92
rect 734 88 738 92
rect 934 88 938 92
rect 1030 88 1034 92
rect 1326 88 1330 92
rect 1366 88 1370 92
rect 1406 88 1410 92
rect 1414 88 1418 92
rect 182 78 186 82
rect 278 78 282 82
rect 334 78 338 82
rect 430 78 434 82
rect 446 78 450 82
rect 486 78 490 82
rect 494 78 498 82
rect 614 78 618 82
rect 646 78 650 82
rect 726 78 730 82
rect 814 78 818 82
rect 918 78 922 82
rect 1038 78 1042 82
rect 1046 78 1050 82
rect 1086 78 1090 82
rect 1126 78 1130 82
rect 1142 78 1146 82
rect 1238 78 1242 82
rect 1334 78 1338 82
rect 1398 79 1402 83
rect 1422 79 1426 83
rect 30 68 34 72
rect 166 68 170 72
rect 302 68 306 72
rect 318 68 322 72
rect 350 68 354 72
rect 422 68 426 72
rect 470 68 474 72
rect 510 68 514 72
rect 526 68 530 72
rect 582 68 586 72
rect 590 68 594 72
rect 606 68 610 72
rect 702 68 706 72
rect 830 68 834 72
rect 942 68 946 72
rect 950 68 954 72
rect 982 68 986 72
rect 1022 68 1026 72
rect 1118 68 1122 72
rect 1254 68 1258 72
rect 6 58 10 62
rect 222 58 226 62
rect 294 58 298 62
rect 326 58 330 62
rect 358 58 362 62
rect 414 58 418 62
rect 462 58 466 62
rect 534 58 538 62
rect 550 58 554 62
rect 574 58 578 62
rect 630 58 634 62
rect 670 58 674 62
rect 694 58 698 62
rect 774 58 778 62
rect 902 58 906 62
rect 958 58 962 62
rect 974 58 978 62
rect 1014 58 1018 62
rect 1070 58 1074 62
rect 1094 58 1098 62
rect 1110 58 1114 62
rect 1126 58 1130 62
rect 1302 58 1306 62
rect 1334 58 1338 62
rect 1390 58 1394 62
rect 1430 58 1434 62
rect 118 48 122 52
rect 390 48 394 52
rect 398 48 402 52
rect 550 48 554 52
rect 582 48 586 52
rect 678 48 682 52
rect 718 48 722 52
rect 878 48 882 52
rect 1086 48 1090 52
rect 1094 48 1098 52
rect 1302 48 1306 52
rect 14 38 18 42
rect 1358 38 1362 42
rect 774 27 778 31
rect 22 18 26 22
rect 118 18 122 22
rect 1302 18 1306 22
rect 442 3 446 7
rect 449 3 453 7
<< metal2 >>
rect 62 1331 66 1332
rect 270 1331 274 1332
rect 62 1328 73 1331
rect 6 1252 9 1268
rect 10 1218 14 1221
rect 30 1192 33 1298
rect 38 1272 41 1288
rect 22 1152 25 1158
rect 46 1152 49 1218
rect 6 1142 9 1148
rect 14 1082 17 1148
rect 54 1142 57 1148
rect 62 1101 65 1258
rect 70 1192 73 1328
rect 262 1328 274 1331
rect 486 1331 490 1332
rect 934 1331 938 1332
rect 486 1328 497 1331
rect 262 1292 265 1328
rect 494 1292 497 1328
rect 926 1328 938 1331
rect 998 1328 1002 1332
rect 1014 1328 1018 1332
rect 1302 1328 1306 1332
rect 1318 1328 1322 1332
rect 1334 1331 1338 1332
rect 1350 1331 1354 1332
rect 1326 1328 1338 1331
rect 1342 1328 1354 1331
rect 1366 1328 1370 1332
rect 1382 1328 1386 1332
rect 1398 1328 1402 1332
rect 1414 1328 1418 1332
rect 1430 1328 1434 1332
rect 926 1292 929 1328
rect 960 1303 962 1307
rect 966 1303 969 1307
rect 973 1303 976 1307
rect 998 1302 1001 1328
rect 1014 1292 1017 1328
rect 1302 1302 1305 1328
rect 1206 1292 1209 1298
rect 1278 1292 1281 1298
rect 1318 1292 1321 1328
rect 1326 1292 1329 1328
rect 1342 1321 1345 1328
rect 1334 1318 1345 1321
rect 1334 1292 1337 1318
rect 1366 1302 1369 1328
rect 978 1288 982 1291
rect 1186 1288 1190 1291
rect 1258 1288 1262 1291
rect 754 1278 758 1281
rect 1166 1279 1174 1281
rect 1190 1279 1198 1281
rect 1214 1279 1222 1281
rect 1230 1282 1233 1288
rect 1166 1278 1177 1279
rect 1190 1278 1201 1279
rect 1214 1278 1225 1279
rect 1238 1279 1246 1281
rect 1262 1279 1270 1281
rect 1286 1279 1294 1281
rect 1302 1282 1305 1288
rect 1238 1278 1249 1279
rect 1262 1278 1273 1279
rect 1286 1278 1297 1279
rect 90 1218 94 1221
rect 174 1221 177 1278
rect 190 1242 193 1268
rect 298 1258 302 1261
rect 166 1218 177 1221
rect 85 1152 88 1158
rect 166 1142 169 1218
rect 182 1152 185 1178
rect 230 1162 233 1258
rect 278 1252 281 1258
rect 238 1222 241 1248
rect 54 1098 65 1101
rect 6 901 9 1018
rect 14 992 17 1078
rect 38 1022 41 1048
rect 6 898 17 901
rect 6 862 9 888
rect 6 761 9 858
rect 14 772 17 898
rect 30 862 33 868
rect 46 862 49 1058
rect 54 952 57 1098
rect 102 1082 105 1138
rect 166 1132 169 1138
rect 182 1132 185 1138
rect 86 1072 89 1078
rect 214 1072 217 1156
rect 254 1142 257 1218
rect 294 1192 297 1238
rect 302 1222 305 1248
rect 350 1192 353 1268
rect 270 1132 273 1158
rect 222 1082 225 1088
rect 270 1072 273 1128
rect 302 1112 305 1138
rect 302 1072 305 1098
rect 310 1092 313 1158
rect 334 1152 337 1158
rect 346 1148 350 1151
rect 326 1072 329 1148
rect 366 1142 369 1278
rect 502 1272 505 1278
rect 518 1262 521 1278
rect 474 1258 478 1261
rect 334 1102 337 1138
rect 342 1122 345 1138
rect 374 1132 377 1158
rect 398 1142 401 1188
rect 406 1152 409 1258
rect 440 1203 442 1207
rect 446 1203 449 1207
rect 453 1203 456 1207
rect 470 1192 473 1238
rect 534 1212 537 1218
rect 446 1160 449 1179
rect 426 1148 430 1151
rect 478 1142 481 1168
rect 534 1162 537 1208
rect 494 1132 497 1138
rect 282 1068 286 1071
rect 142 1062 145 1068
rect 238 1062 241 1068
rect 214 1052 217 1058
rect 194 1048 198 1051
rect 246 1042 249 1068
rect 270 1062 273 1068
rect 294 1062 297 1068
rect 282 1058 286 1061
rect 302 1032 305 1068
rect 334 1062 337 1088
rect 342 1062 345 1068
rect 310 1052 313 1058
rect 334 1052 337 1058
rect 358 1052 361 1128
rect 366 992 369 1118
rect 494 1111 497 1128
rect 494 1108 505 1111
rect 502 1082 505 1108
rect 502 1072 505 1078
rect 378 1068 382 1071
rect 382 1052 385 1058
rect 398 1051 401 1068
rect 410 1058 414 1061
rect 518 1052 521 1068
rect 574 1062 577 1258
rect 582 1152 585 1158
rect 590 1142 593 1208
rect 606 1132 609 1158
rect 398 1048 409 1051
rect 390 992 393 1038
rect 158 962 161 988
rect 198 962 201 988
rect 166 952 169 958
rect 302 952 305 958
rect 194 948 198 951
rect 378 948 382 951
rect 110 932 113 938
rect 94 912 97 928
rect 118 882 121 908
rect 102 872 105 878
rect 50 858 54 861
rect 54 822 57 848
rect 62 792 65 848
rect 102 792 105 858
rect 118 852 121 878
rect 110 772 113 808
rect 158 792 161 868
rect 198 772 201 948
rect 218 878 222 881
rect 230 872 233 878
rect 246 872 249 938
rect 346 928 350 931
rect 378 928 382 931
rect 262 912 265 928
rect 262 882 265 908
rect 6 758 17 761
rect 6 722 9 738
rect 6 492 9 718
rect 14 712 17 758
rect 86 752 89 758
rect 110 752 113 768
rect 222 762 225 818
rect 130 758 134 761
rect 150 752 153 758
rect 122 748 126 751
rect 14 481 17 708
rect 134 692 137 728
rect 162 688 166 691
rect 174 682 177 748
rect 70 672 73 678
rect 22 622 25 648
rect 22 562 25 588
rect 38 552 41 658
rect 6 478 17 481
rect 22 492 25 548
rect 70 542 73 548
rect 86 532 89 678
rect 182 642 185 748
rect 190 682 193 728
rect 222 692 225 758
rect 238 752 241 758
rect 246 752 249 798
rect 262 752 265 878
rect 278 862 281 868
rect 286 862 289 908
rect 302 882 305 918
rect 318 892 321 928
rect 338 918 342 921
rect 298 858 302 861
rect 286 802 289 858
rect 310 812 313 878
rect 334 872 337 898
rect 358 892 361 928
rect 398 882 401 1038
rect 406 992 409 1048
rect 410 948 414 951
rect 422 942 425 948
rect 430 942 433 1028
rect 440 1003 442 1007
rect 446 1003 449 1007
rect 453 1003 456 1007
rect 478 992 481 1008
rect 438 982 441 988
rect 482 948 486 951
rect 522 948 526 951
rect 494 942 497 948
rect 514 938 518 941
rect 342 862 345 868
rect 358 842 361 848
rect 270 752 273 768
rect 286 760 289 779
rect 390 762 393 838
rect 398 792 401 878
rect 406 802 409 818
rect 410 788 414 791
rect 422 782 425 928
rect 462 921 465 928
rect 494 922 497 938
rect 534 932 537 968
rect 462 918 470 921
rect 390 752 393 758
rect 230 732 233 738
rect 318 732 321 738
rect 334 732 337 748
rect 430 742 433 898
rect 486 882 489 888
rect 502 862 505 868
rect 550 862 553 1058
rect 574 1052 577 1058
rect 582 1051 585 1088
rect 614 1072 617 1278
rect 734 1272 737 1278
rect 630 1192 633 1268
rect 702 1262 705 1268
rect 682 1258 686 1261
rect 722 1258 726 1261
rect 678 1222 681 1248
rect 798 1231 801 1258
rect 718 1162 721 1168
rect 630 1138 638 1141
rect 622 1072 625 1138
rect 630 1092 633 1138
rect 646 1092 649 1158
rect 666 1148 670 1151
rect 674 1138 678 1141
rect 694 1132 697 1158
rect 726 1152 729 1158
rect 734 1152 737 1188
rect 742 1182 745 1218
rect 782 1162 785 1168
rect 758 1152 761 1158
rect 790 1152 793 1158
rect 770 1148 774 1151
rect 802 1148 806 1151
rect 694 1112 697 1128
rect 590 1062 593 1068
rect 610 1058 614 1061
rect 582 1048 590 1051
rect 566 1022 569 1048
rect 622 992 625 1058
rect 638 1012 641 1078
rect 646 1062 649 1078
rect 670 1062 673 1088
rect 690 1078 694 1081
rect 710 1062 713 1148
rect 786 1138 790 1141
rect 726 1082 729 1138
rect 706 1058 710 1061
rect 646 1042 649 1058
rect 702 1032 705 1038
rect 718 1002 721 1048
rect 726 991 729 1058
rect 734 1032 737 1138
rect 798 1132 801 1138
rect 822 1132 825 1138
rect 758 1092 761 1128
rect 830 1112 833 1158
rect 838 1102 841 1278
rect 1078 1272 1081 1278
rect 854 1212 857 1268
rect 906 1248 910 1251
rect 942 1222 945 1258
rect 870 1192 873 1208
rect 846 1152 849 1158
rect 854 1152 857 1158
rect 862 1152 865 1178
rect 846 1142 849 1148
rect 862 1082 865 1118
rect 746 1078 750 1081
rect 766 1062 769 1078
rect 746 1058 750 1061
rect 778 1038 782 1041
rect 722 988 729 991
rect 790 992 793 1078
rect 862 1072 865 1078
rect 878 1072 881 1078
rect 822 1052 825 1058
rect 830 992 833 1008
rect 862 992 865 1058
rect 910 1031 913 1050
rect 566 962 569 978
rect 562 958 566 961
rect 606 952 609 978
rect 706 968 710 971
rect 718 952 721 988
rect 838 972 841 988
rect 910 972 913 1008
rect 918 992 921 1148
rect 925 1142 928 1148
rect 934 1062 937 1148
rect 950 1092 953 1258
rect 1038 1252 1041 1258
rect 1002 1218 1006 1221
rect 1094 1221 1097 1268
rect 1166 1262 1169 1278
rect 1190 1262 1193 1278
rect 1214 1262 1217 1278
rect 1238 1262 1241 1278
rect 1086 1218 1097 1221
rect 1054 1160 1057 1179
rect 962 1148 966 1151
rect 1022 1132 1025 1138
rect 1006 1122 1009 1128
rect 960 1103 962 1107
rect 966 1103 969 1107
rect 973 1103 976 1107
rect 1006 1092 1009 1108
rect 1030 1092 1033 1108
rect 966 1072 969 1088
rect 1050 1078 1054 1081
rect 950 1052 953 1068
rect 1010 1058 1014 1061
rect 962 1048 966 1051
rect 874 968 894 971
rect 850 958 854 961
rect 726 952 729 958
rect 802 948 806 951
rect 742 942 745 948
rect 606 932 609 938
rect 738 928 742 931
rect 622 912 625 928
rect 654 882 657 908
rect 750 902 753 948
rect 766 942 769 948
rect 758 932 761 938
rect 738 888 742 891
rect 534 831 537 850
rect 440 803 442 807
rect 446 803 449 807
rect 453 803 456 807
rect 478 792 481 818
rect 558 792 561 868
rect 586 858 590 861
rect 438 772 441 778
rect 458 758 462 761
rect 438 752 441 758
rect 486 702 489 728
rect 422 692 425 698
rect 502 692 505 718
rect 518 712 521 748
rect 526 732 529 788
rect 574 752 577 758
rect 198 682 201 688
rect 170 588 174 591
rect 182 552 185 618
rect 190 592 193 678
rect 218 668 222 671
rect 246 662 249 688
rect 342 682 345 688
rect 518 682 521 698
rect 534 682 537 718
rect 450 678 454 681
rect 254 642 257 658
rect 214 552 217 618
rect 222 552 225 638
rect 278 622 281 648
rect 246 562 249 588
rect 294 552 297 658
rect 326 652 329 668
rect 390 592 393 678
rect 502 662 505 668
rect 510 662 513 668
rect 518 662 521 668
rect 566 662 569 678
rect 574 662 577 668
rect 582 662 585 748
rect 590 722 593 738
rect 598 682 601 878
rect 606 831 609 850
rect 638 812 641 868
rect 654 821 657 878
rect 646 818 657 821
rect 646 792 649 818
rect 678 792 681 808
rect 710 762 713 768
rect 670 752 673 758
rect 706 748 710 751
rect 598 672 601 678
rect 606 672 609 748
rect 694 742 697 748
rect 718 732 721 888
rect 774 872 777 938
rect 782 902 785 948
rect 782 892 785 898
rect 790 882 793 948
rect 814 932 817 938
rect 806 892 809 898
rect 798 872 801 878
rect 734 762 737 848
rect 742 792 745 838
rect 750 782 753 868
rect 814 852 817 858
rect 762 848 766 851
rect 822 842 825 958
rect 858 948 862 951
rect 774 792 777 838
rect 830 792 833 948
rect 862 892 865 918
rect 886 902 889 958
rect 910 942 913 968
rect 950 962 953 1048
rect 966 952 969 1018
rect 990 1012 993 1058
rect 1022 1022 1025 1068
rect 1062 1062 1065 1098
rect 1070 1082 1073 1218
rect 1086 1112 1089 1218
rect 1134 1212 1137 1258
rect 1142 1222 1145 1248
rect 1130 1138 1134 1141
rect 1094 1081 1097 1128
rect 1118 1102 1121 1138
rect 1142 1102 1145 1148
rect 1158 1092 1161 1128
rect 1086 1078 1097 1081
rect 1070 1062 1073 1078
rect 1078 1062 1081 1068
rect 1062 1022 1065 1058
rect 1086 1032 1089 1078
rect 1154 1068 1158 1071
rect 1094 1032 1097 1068
rect 1102 1052 1105 1058
rect 986 988 990 991
rect 1030 952 1033 1008
rect 1038 992 1041 998
rect 1050 968 1054 971
rect 1086 962 1089 978
rect 1094 972 1097 1018
rect 1110 1012 1113 1068
rect 1118 1062 1121 1068
rect 1122 1048 1126 1051
rect 1134 992 1137 1068
rect 1190 1062 1193 1208
rect 1254 1132 1257 1268
rect 1262 1262 1265 1278
rect 1286 1262 1289 1278
rect 1310 1241 1313 1258
rect 1310 1238 1318 1241
rect 1334 1202 1337 1258
rect 1350 1251 1353 1298
rect 1374 1292 1377 1298
rect 1382 1292 1385 1328
rect 1398 1302 1401 1328
rect 1414 1302 1417 1328
rect 1430 1302 1433 1328
rect 1358 1279 1366 1281
rect 1382 1279 1390 1281
rect 1406 1279 1414 1281
rect 1358 1278 1369 1279
rect 1382 1278 1393 1279
rect 1406 1278 1417 1279
rect 1358 1262 1361 1278
rect 1382 1262 1385 1278
rect 1406 1262 1409 1278
rect 1350 1248 1361 1251
rect 1350 1222 1353 1228
rect 1358 1192 1361 1248
rect 1270 1152 1273 1178
rect 1270 1132 1273 1138
rect 1254 1101 1257 1128
rect 1246 1098 1257 1101
rect 1246 1082 1249 1098
rect 1302 1092 1305 1156
rect 1230 1072 1233 1078
rect 1286 1062 1289 1088
rect 1342 1062 1345 1148
rect 1358 1092 1361 1168
rect 1366 1152 1369 1208
rect 1390 1152 1393 1208
rect 1398 1182 1401 1218
rect 1414 1152 1417 1208
rect 1406 1132 1409 1138
rect 1422 1122 1425 1278
rect 1434 1238 1438 1241
rect 1382 1102 1385 1118
rect 1406 1092 1409 1118
rect 1366 1079 1374 1081
rect 1366 1078 1377 1079
rect 1366 1062 1369 1078
rect 1438 1062 1441 1118
rect 1158 1052 1161 1058
rect 1190 982 1193 1058
rect 1198 1031 1201 1050
rect 1230 992 1233 1058
rect 1382 1022 1385 1028
rect 1326 1012 1329 1018
rect 1390 992 1393 1058
rect 1414 1002 1417 1058
rect 1438 1032 1441 1038
rect 1438 992 1441 1008
rect 1402 988 1406 991
rect 954 948 958 951
rect 1010 948 1014 951
rect 1050 948 1054 951
rect 950 932 953 938
rect 958 932 961 948
rect 910 912 913 928
rect 966 922 969 948
rect 960 903 962 907
rect 966 903 969 907
rect 973 903 976 907
rect 914 888 918 891
rect 862 862 865 868
rect 850 858 854 861
rect 862 792 865 848
rect 870 842 873 878
rect 730 758 734 761
rect 742 752 745 778
rect 770 768 774 771
rect 826 768 830 771
rect 774 742 777 748
rect 750 722 753 738
rect 782 722 785 758
rect 830 752 833 758
rect 794 748 798 751
rect 686 662 689 688
rect 726 682 729 688
rect 742 672 745 678
rect 578 658 582 661
rect 510 642 513 658
rect 550 652 553 658
rect 438 622 441 628
rect 440 603 442 607
rect 446 603 449 607
rect 453 603 456 607
rect 178 538 182 541
rect 246 532 249 548
rect 486 542 489 618
rect 590 602 593 618
rect 494 562 497 588
rect 606 562 609 658
rect 614 612 617 618
rect 638 592 641 638
rect 646 582 649 618
rect 502 552 505 558
rect 542 542 545 548
rect 294 532 297 538
rect 86 522 89 528
rect 6 462 9 478
rect 22 462 25 488
rect 118 482 121 508
rect 102 472 105 478
rect 158 462 161 468
rect 230 462 233 528
rect 310 512 313 528
rect 294 482 297 508
rect 278 462 281 468
rect 50 458 54 461
rect 226 458 230 461
rect 6 352 9 458
rect 54 422 57 448
rect 202 428 206 431
rect 246 431 249 450
rect 54 362 57 388
rect 246 360 249 379
rect 206 352 209 358
rect 50 348 54 351
rect 226 348 230 351
rect 22 322 25 348
rect 102 332 105 338
rect 22 262 25 318
rect 118 312 121 328
rect 86 282 89 308
rect 70 262 73 268
rect 22 222 25 248
rect 62 192 65 218
rect 10 138 14 141
rect 30 72 33 138
rect 86 132 89 278
rect 126 262 129 268
rect 198 262 201 348
rect 278 342 281 348
rect 294 332 297 478
rect 398 472 401 538
rect 422 482 425 518
rect 438 492 441 532
rect 558 522 561 528
rect 446 482 449 508
rect 410 458 414 461
rect 378 448 382 451
rect 374 392 377 438
rect 390 432 393 448
rect 422 422 425 458
rect 294 312 297 328
rect 262 282 265 308
rect 246 272 249 278
rect 194 258 198 261
rect 170 238 174 241
rect 190 201 193 258
rect 198 222 201 248
rect 262 222 265 278
rect 190 198 201 201
rect 94 162 97 188
rect 198 152 201 198
rect 238 162 241 168
rect 142 142 145 148
rect 86 92 89 128
rect 158 122 161 128
rect 158 102 161 118
rect 198 102 201 148
rect 294 122 297 148
rect 302 132 305 248
rect 310 142 313 158
rect 318 142 321 188
rect 334 162 337 348
rect 398 342 401 358
rect 422 352 425 358
rect 430 341 433 468
rect 470 462 473 468
rect 478 462 481 498
rect 590 492 593 498
rect 526 482 529 488
rect 598 482 601 498
rect 554 478 558 481
rect 610 478 614 481
rect 486 462 489 468
rect 494 462 497 468
rect 440 403 442 407
rect 446 403 449 407
rect 453 403 456 407
rect 470 372 473 458
rect 430 338 438 341
rect 442 338 446 341
rect 390 302 393 318
rect 390 282 393 298
rect 398 272 401 278
rect 374 262 377 268
rect 406 262 409 288
rect 418 268 422 271
rect 418 258 422 261
rect 430 261 433 328
rect 438 272 441 308
rect 454 282 457 338
rect 470 282 473 368
rect 478 352 481 418
rect 502 412 505 468
rect 518 452 521 468
rect 526 462 529 478
rect 550 462 553 478
rect 630 462 633 578
rect 658 568 662 571
rect 686 552 689 578
rect 694 562 697 568
rect 702 562 705 608
rect 726 552 729 638
rect 774 631 777 650
rect 782 632 785 658
rect 790 582 793 748
rect 798 732 801 738
rect 806 732 809 738
rect 798 682 801 728
rect 814 692 817 698
rect 838 691 841 748
rect 854 702 857 768
rect 870 762 873 768
rect 878 762 881 878
rect 942 872 945 878
rect 922 858 926 861
rect 886 792 889 858
rect 902 852 905 858
rect 862 752 865 758
rect 878 742 881 758
rect 886 752 889 768
rect 838 688 849 691
rect 834 678 838 681
rect 830 662 833 668
rect 734 562 737 568
rect 774 552 777 558
rect 798 552 801 658
rect 818 648 822 651
rect 830 562 833 618
rect 846 562 849 688
rect 854 662 857 668
rect 870 662 873 718
rect 894 712 897 768
rect 910 742 913 748
rect 918 711 921 848
rect 930 768 934 771
rect 942 752 945 868
rect 970 858 974 861
rect 966 792 969 818
rect 966 752 969 758
rect 942 732 945 748
rect 914 708 921 711
rect 886 692 889 698
rect 910 692 913 708
rect 926 692 929 718
rect 950 692 953 728
rect 960 703 962 707
rect 966 703 969 707
rect 973 703 976 707
rect 982 702 985 878
rect 998 772 1001 928
rect 1006 892 1009 928
rect 1022 912 1025 938
rect 1062 922 1065 958
rect 1134 952 1137 978
rect 1262 952 1265 978
rect 1278 960 1281 979
rect 1134 932 1137 938
rect 1150 932 1153 938
rect 1014 882 1017 888
rect 1042 878 1046 881
rect 1006 872 1009 878
rect 1026 868 1030 871
rect 1006 852 1009 858
rect 1046 852 1049 868
rect 1054 862 1057 868
rect 990 742 993 748
rect 998 692 1001 748
rect 1006 722 1009 848
rect 1054 752 1057 858
rect 1070 792 1073 908
rect 1134 892 1137 918
rect 1122 888 1126 891
rect 1162 878 1166 881
rect 1082 858 1086 861
rect 1106 858 1110 861
rect 1118 852 1121 868
rect 1078 781 1081 848
rect 1126 842 1129 878
rect 1174 872 1177 878
rect 1190 872 1193 938
rect 1226 918 1230 921
rect 1202 868 1206 871
rect 1166 862 1169 868
rect 1230 862 1233 888
rect 1242 868 1246 871
rect 1262 862 1265 948
rect 1310 942 1313 948
rect 1326 882 1329 928
rect 1110 792 1113 838
rect 1142 832 1145 848
rect 1074 778 1081 781
rect 1022 692 1025 728
rect 1030 692 1033 728
rect 1046 722 1049 748
rect 1070 692 1073 778
rect 1126 771 1129 828
rect 1142 792 1145 818
rect 1174 772 1177 828
rect 1182 822 1185 848
rect 1182 792 1185 808
rect 1126 768 1134 771
rect 1094 752 1097 758
rect 1086 742 1089 748
rect 1102 732 1105 758
rect 1114 738 1118 741
rect 1126 692 1129 768
rect 1150 762 1153 768
rect 1142 742 1145 748
rect 1166 742 1169 748
rect 1118 682 1121 688
rect 946 678 950 681
rect 1042 678 1046 681
rect 894 672 897 678
rect 878 662 881 668
rect 902 662 905 678
rect 918 662 921 678
rect 930 668 934 671
rect 858 648 862 651
rect 854 562 857 588
rect 786 548 790 551
rect 658 528 665 531
rect 662 502 665 528
rect 662 492 665 498
rect 670 492 673 538
rect 678 492 681 548
rect 702 542 705 548
rect 786 538 790 541
rect 750 532 753 538
rect 646 472 649 478
rect 578 458 582 461
rect 566 452 569 458
rect 518 402 521 448
rect 430 258 438 261
rect 454 252 457 278
rect 478 272 481 348
rect 486 342 489 358
rect 510 332 513 348
rect 526 342 529 388
rect 534 332 537 418
rect 566 392 569 448
rect 566 362 569 368
rect 574 362 577 378
rect 582 362 585 418
rect 598 392 601 458
rect 622 432 625 458
rect 630 452 633 458
rect 638 441 641 468
rect 634 438 641 441
rect 654 442 657 478
rect 678 472 681 478
rect 670 462 673 468
rect 678 462 681 468
rect 654 422 657 438
rect 542 358 550 361
rect 498 328 502 331
rect 514 328 518 331
rect 494 312 497 318
rect 542 302 545 358
rect 606 352 609 398
rect 654 362 657 398
rect 614 352 617 358
rect 570 348 574 351
rect 550 342 553 348
rect 626 338 630 341
rect 626 328 630 331
rect 590 322 593 328
rect 494 282 497 288
rect 478 252 481 258
rect 342 222 345 228
rect 374 192 377 218
rect 440 203 442 207
rect 446 203 449 207
rect 453 203 456 207
rect 334 142 337 158
rect 350 152 353 188
rect 366 172 369 178
rect 398 162 401 178
rect 378 148 382 151
rect 394 148 398 151
rect 422 142 425 158
rect 438 142 441 168
rect 446 152 449 188
rect 478 152 481 158
rect 502 152 505 278
rect 510 272 513 278
rect 510 182 513 268
rect 526 262 529 298
rect 546 268 550 271
rect 558 262 561 318
rect 598 282 601 288
rect 606 272 609 278
rect 578 268 582 271
rect 538 238 542 241
rect 510 162 513 168
rect 458 148 462 151
rect 490 138 494 141
rect 374 122 377 138
rect 406 132 409 138
rect 418 128 422 131
rect 430 122 433 128
rect 182 82 185 98
rect 166 72 169 78
rect 222 62 225 98
rect 282 78 286 81
rect 318 72 321 88
rect 298 68 302 71
rect 326 62 329 98
rect 334 82 337 118
rect 394 88 398 91
rect 350 72 353 78
rect 422 72 425 88
rect 450 78 454 81
rect 430 72 433 78
rect 354 68 358 71
rect 462 62 465 138
rect 478 132 481 138
rect 494 122 497 138
rect 502 92 505 98
rect 482 88 486 91
rect 482 78 486 81
rect 486 72 489 78
rect 470 62 473 68
rect 298 58 302 61
rect 362 58 366 61
rect 410 58 414 61
rect 6 41 9 58
rect 390 52 393 58
rect 494 52 497 78
rect 510 72 513 158
rect 534 152 537 198
rect 542 142 545 228
rect 558 222 561 258
rect 574 242 577 248
rect 582 232 585 258
rect 590 242 593 248
rect 550 132 553 138
rect 558 132 561 178
rect 566 162 569 228
rect 614 152 617 288
rect 622 282 625 318
rect 638 301 641 338
rect 634 298 641 301
rect 630 272 633 298
rect 646 282 649 348
rect 678 342 681 348
rect 670 321 673 338
rect 686 331 689 528
rect 750 492 753 518
rect 758 482 761 538
rect 778 528 785 531
rect 774 512 777 518
rect 774 502 777 508
rect 782 492 785 528
rect 798 492 801 538
rect 806 492 809 558
rect 862 552 865 628
rect 774 472 777 488
rect 798 482 801 488
rect 790 472 793 478
rect 814 472 817 538
rect 870 532 873 658
rect 926 622 929 668
rect 990 662 993 678
rect 1014 672 1017 678
rect 1078 672 1081 678
rect 1002 668 1006 671
rect 1014 652 1017 668
rect 1046 662 1049 668
rect 1078 662 1081 668
rect 1134 662 1137 718
rect 1174 712 1177 768
rect 1190 732 1193 838
rect 1198 832 1201 858
rect 1310 852 1313 868
rect 1214 812 1217 848
rect 1230 842 1233 848
rect 1278 831 1281 850
rect 1238 792 1241 828
rect 1326 812 1329 878
rect 1414 862 1417 888
rect 1422 862 1425 948
rect 1438 892 1441 968
rect 1402 858 1407 861
rect 1210 748 1214 751
rect 1206 722 1209 738
rect 1342 732 1345 808
rect 1390 760 1393 779
rect 1062 652 1065 658
rect 1098 648 1102 651
rect 934 642 937 648
rect 902 542 905 548
rect 918 532 921 598
rect 998 592 1001 598
rect 1010 538 1014 541
rect 1034 528 1038 531
rect 830 512 833 518
rect 960 503 962 507
rect 966 503 969 507
rect 973 503 976 507
rect 754 468 758 471
rect 694 452 697 458
rect 702 452 705 468
rect 726 452 729 468
rect 694 432 697 448
rect 694 342 697 398
rect 702 382 705 448
rect 710 392 713 418
rect 726 402 729 448
rect 734 432 737 468
rect 822 462 825 468
rect 830 462 833 468
rect 838 462 841 498
rect 874 488 878 491
rect 902 472 905 498
rect 918 472 921 478
rect 882 468 886 471
rect 926 462 929 498
rect 962 488 966 491
rect 934 472 937 478
rect 882 458 886 461
rect 914 458 918 461
rect 766 452 769 458
rect 746 448 750 451
rect 734 352 737 408
rect 758 372 761 428
rect 706 348 710 351
rect 742 342 745 358
rect 758 351 761 368
rect 766 362 769 368
rect 774 352 777 388
rect 794 368 798 371
rect 806 362 809 448
rect 786 358 790 361
rect 758 348 769 351
rect 794 348 809 351
rect 682 328 689 331
rect 706 328 710 331
rect 670 318 681 321
rect 630 252 633 258
rect 630 192 633 228
rect 638 202 641 258
rect 646 252 649 258
rect 654 252 657 318
rect 678 292 681 318
rect 666 258 673 261
rect 662 192 665 198
rect 670 152 673 258
rect 686 222 689 328
rect 694 272 697 308
rect 718 281 721 318
rect 726 302 729 328
rect 742 292 745 338
rect 750 302 753 348
rect 766 292 769 348
rect 774 322 777 328
rect 782 312 785 348
rect 718 278 729 281
rect 726 272 729 278
rect 714 268 718 271
rect 702 242 705 258
rect 738 248 742 251
rect 686 182 689 218
rect 718 181 721 248
rect 726 192 729 218
rect 734 192 737 248
rect 718 178 729 181
rect 602 148 606 151
rect 650 148 654 151
rect 674 148 678 151
rect 714 148 718 151
rect 638 142 641 148
rect 586 138 590 141
rect 614 122 617 138
rect 518 82 521 118
rect 554 88 558 91
rect 522 68 526 71
rect 402 48 406 51
rect 6 38 14 41
rect 118 22 121 48
rect 534 42 537 58
rect 542 51 545 78
rect 582 72 585 98
rect 614 82 617 118
rect 622 92 625 128
rect 646 82 649 88
rect 590 72 593 78
rect 574 62 577 68
rect 554 58 558 61
rect 582 52 585 68
rect 606 62 609 68
rect 634 58 638 61
rect 542 48 550 51
rect 646 42 649 78
rect 670 62 673 148
rect 698 138 702 141
rect 726 82 729 178
rect 738 148 742 151
rect 750 151 753 258
rect 758 192 761 278
rect 782 272 785 308
rect 790 292 793 338
rect 798 312 801 338
rect 806 322 809 348
rect 814 342 817 398
rect 822 362 825 458
rect 894 452 897 458
rect 858 448 862 451
rect 874 358 878 361
rect 822 342 825 348
rect 846 342 849 358
rect 878 342 881 348
rect 886 342 889 398
rect 926 392 929 448
rect 918 362 921 368
rect 902 352 905 358
rect 826 328 830 331
rect 806 272 809 298
rect 822 292 825 298
rect 830 282 833 318
rect 838 312 841 318
rect 862 302 865 338
rect 886 272 889 298
rect 866 268 870 271
rect 798 232 801 248
rect 746 148 753 151
rect 734 92 737 148
rect 798 141 801 198
rect 806 152 809 268
rect 822 252 825 258
rect 830 152 833 238
rect 798 138 806 141
rect 814 132 817 148
rect 838 101 841 248
rect 846 222 849 268
rect 878 262 881 268
rect 854 202 857 258
rect 862 191 865 248
rect 858 188 865 191
rect 878 192 881 228
rect 830 98 841 101
rect 858 148 862 151
rect 854 102 857 148
rect 862 132 865 138
rect 878 131 881 148
rect 886 132 889 268
rect 894 212 897 348
rect 910 342 913 358
rect 902 272 905 328
rect 934 312 937 338
rect 942 331 945 478
rect 1006 472 1009 478
rect 954 468 958 471
rect 950 342 953 468
rect 1006 462 1009 468
rect 1022 462 1025 488
rect 1046 482 1049 488
rect 966 372 969 448
rect 974 352 977 388
rect 942 328 953 331
rect 942 302 945 318
rect 930 278 934 281
rect 902 242 905 268
rect 910 232 913 258
rect 894 142 897 148
rect 902 142 905 218
rect 910 162 913 218
rect 926 202 929 278
rect 950 262 953 328
rect 960 303 962 307
rect 966 303 969 307
rect 973 303 976 307
rect 982 292 985 458
rect 998 452 1001 458
rect 1006 362 1009 458
rect 1030 442 1033 478
rect 1054 472 1057 558
rect 1070 552 1073 588
rect 1062 462 1065 548
rect 1078 542 1081 578
rect 1110 562 1113 568
rect 1150 552 1153 558
rect 1158 552 1161 618
rect 1174 592 1177 698
rect 1190 692 1193 708
rect 1182 682 1185 688
rect 1186 668 1190 671
rect 1198 662 1201 718
rect 1242 618 1246 621
rect 1262 602 1265 718
rect 1342 712 1345 728
rect 1358 712 1361 738
rect 1326 682 1329 708
rect 1286 632 1289 658
rect 1238 552 1241 598
rect 1286 591 1289 628
rect 1286 588 1297 591
rect 1294 552 1297 588
rect 1106 548 1110 551
rect 1110 522 1113 538
rect 1086 482 1089 518
rect 1094 482 1097 518
rect 1058 438 1062 441
rect 1074 438 1078 441
rect 1086 432 1089 458
rect 1094 452 1097 478
rect 1102 442 1105 478
rect 1118 472 1121 548
rect 1134 542 1137 548
rect 1134 532 1137 538
rect 1150 532 1153 538
rect 1134 491 1137 528
rect 1158 522 1161 548
rect 1194 538 1197 541
rect 1190 502 1193 528
rect 1130 488 1137 491
rect 1126 462 1129 488
rect 1198 482 1201 538
rect 1218 488 1222 491
rect 1138 478 1142 481
rect 1170 478 1174 481
rect 1150 472 1153 478
rect 1238 472 1241 548
rect 1278 532 1281 538
rect 1294 511 1297 538
rect 1326 532 1329 678
rect 1342 621 1345 668
rect 1374 631 1377 650
rect 1334 618 1345 621
rect 1286 508 1297 511
rect 1286 492 1289 508
rect 1258 488 1265 491
rect 1262 482 1265 488
rect 1250 478 1254 481
rect 1274 478 1278 481
rect 1294 472 1297 488
rect 1326 482 1329 518
rect 1334 482 1337 618
rect 1342 562 1345 588
rect 1366 532 1369 538
rect 1382 492 1385 708
rect 1398 662 1401 748
rect 1414 611 1417 658
rect 1438 642 1441 648
rect 1414 608 1425 611
rect 1350 472 1353 478
rect 1406 472 1409 478
rect 1138 468 1142 471
rect 1162 468 1166 471
rect 1178 468 1182 471
rect 1258 468 1262 471
rect 1166 452 1169 458
rect 1190 452 1193 468
rect 1222 462 1225 468
rect 1238 462 1241 468
rect 1266 458 1270 461
rect 1014 372 1017 378
rect 974 272 977 278
rect 990 262 993 318
rect 1006 272 1009 358
rect 1014 352 1017 358
rect 1022 342 1025 368
rect 1038 342 1041 418
rect 1062 352 1065 358
rect 1046 342 1049 348
rect 1014 338 1022 341
rect 1014 282 1017 338
rect 1038 322 1041 338
rect 1062 332 1065 348
rect 1070 342 1073 348
rect 1078 342 1081 428
rect 1086 362 1089 418
rect 1102 352 1105 418
rect 1126 392 1129 438
rect 1118 342 1121 388
rect 1142 342 1145 368
rect 1154 358 1158 361
rect 1182 352 1185 358
rect 1190 352 1193 358
rect 1198 342 1201 458
rect 1230 452 1233 458
rect 1218 448 1222 451
rect 1302 442 1305 458
rect 1358 452 1361 468
rect 1414 462 1417 558
rect 1406 458 1414 461
rect 1234 368 1238 371
rect 1382 362 1385 388
rect 1406 362 1409 458
rect 1274 348 1278 351
rect 1402 348 1406 351
rect 1206 342 1209 348
rect 1106 338 1110 341
rect 946 258 950 261
rect 958 202 961 238
rect 926 182 929 198
rect 926 152 929 178
rect 966 162 969 168
rect 982 162 985 218
rect 954 158 958 161
rect 914 148 918 151
rect 934 142 937 158
rect 946 148 950 151
rect 922 138 926 141
rect 938 138 945 141
rect 878 128 886 131
rect 914 128 918 131
rect 702 72 705 78
rect 734 72 737 88
rect 814 82 817 88
rect 830 72 833 98
rect 934 92 937 128
rect 922 78 926 81
rect 942 81 945 138
rect 950 91 953 148
rect 966 142 969 148
rect 960 103 962 107
rect 966 103 969 107
rect 973 103 976 107
rect 950 88 961 91
rect 958 82 961 88
rect 942 78 953 81
rect 950 72 953 78
rect 694 62 697 68
rect 718 52 721 58
rect 682 48 686 51
rect 774 31 777 58
rect 878 52 881 68
rect 906 58 910 61
rect 942 52 945 68
rect 950 62 953 68
rect 958 62 961 78
rect 990 72 993 258
rect 1006 222 1009 248
rect 1014 152 1017 198
rect 1014 142 1017 148
rect 974 52 977 58
rect 982 52 985 68
rect 1014 62 1017 128
rect 1022 72 1025 208
rect 1030 192 1033 218
rect 1030 142 1033 148
rect 1030 92 1033 118
rect 1038 82 1041 308
rect 1046 252 1049 318
rect 1102 282 1105 318
rect 1118 282 1121 338
rect 1174 332 1177 338
rect 1222 332 1225 338
rect 1130 328 1134 331
rect 1058 258 1062 261
rect 1102 242 1105 268
rect 1118 262 1121 268
rect 1174 262 1177 268
rect 1054 162 1057 228
rect 1074 158 1081 161
rect 1078 152 1081 158
rect 1066 148 1070 151
rect 1046 132 1049 138
rect 1054 81 1057 138
rect 1050 78 1057 81
rect 1070 62 1073 148
rect 1078 132 1081 138
rect 1102 132 1105 238
rect 1150 231 1153 250
rect 1118 152 1121 178
rect 1134 162 1137 198
rect 1182 192 1185 258
rect 1198 182 1201 218
rect 1214 182 1217 318
rect 1238 272 1241 348
rect 1334 332 1337 338
rect 1318 322 1321 328
rect 1278 282 1281 318
rect 1374 292 1377 318
rect 1238 262 1241 268
rect 1294 262 1297 268
rect 1238 202 1241 258
rect 1342 222 1345 248
rect 1374 202 1377 218
rect 1238 182 1241 188
rect 1202 178 1209 181
rect 1126 152 1129 158
rect 1150 152 1153 178
rect 1198 162 1201 168
rect 1182 152 1185 158
rect 1206 142 1209 178
rect 1214 162 1217 168
rect 1230 162 1233 178
rect 1302 152 1305 198
rect 1258 148 1261 151
rect 1214 142 1217 148
rect 1110 132 1113 138
rect 1078 102 1081 128
rect 1086 82 1089 88
rect 1118 72 1121 78
rect 1126 72 1129 78
rect 1086 52 1089 68
rect 1110 62 1113 68
rect 1098 58 1102 61
rect 1134 61 1137 138
rect 1142 132 1145 138
rect 1254 122 1257 128
rect 1142 82 1145 98
rect 1238 82 1241 108
rect 1130 58 1137 61
rect 1254 62 1257 68
rect 1302 62 1305 148
rect 1342 132 1345 198
rect 1390 160 1393 179
rect 1358 142 1361 148
rect 1342 112 1345 128
rect 1326 92 1329 98
rect 1366 92 1369 108
rect 1406 92 1409 338
rect 1414 92 1417 448
rect 1422 122 1425 608
rect 1430 542 1433 608
rect 1430 272 1433 538
rect 1438 442 1441 448
rect 1438 342 1441 348
rect 1334 82 1337 88
rect 1390 79 1398 81
rect 1426 79 1433 81
rect 1390 78 1401 79
rect 1422 78 1433 79
rect 1390 62 1393 78
rect 1430 62 1433 78
rect 1094 42 1097 48
rect 1302 22 1305 48
rect 14 -19 18 -18
rect 22 -19 25 18
rect 1334 12 1337 58
rect 1358 42 1361 48
rect 440 3 442 7
rect 446 3 449 7
rect 453 3 456 7
rect 14 -22 25 -19
rect 1310 -18 1313 8
rect 1406 -18 1409 8
rect 1422 -18 1425 8
rect 1438 -18 1441 118
rect 1310 -22 1314 -18
rect 1406 -22 1410 -18
rect 1422 -22 1426 -18
rect 1438 -22 1442 -18
<< m3contact >>
rect 30 1298 34 1302
rect 6 1248 10 1252
rect 6 1218 10 1222
rect 38 1288 42 1292
rect 46 1218 50 1222
rect 22 1158 26 1162
rect 6 1148 10 1152
rect 14 1148 18 1152
rect 54 1138 58 1142
rect 962 1303 966 1307
rect 969 1303 973 1307
rect 998 1298 1002 1302
rect 1206 1298 1210 1302
rect 1278 1298 1282 1302
rect 1302 1298 1306 1302
rect 1350 1298 1354 1302
rect 1366 1298 1370 1302
rect 1374 1298 1378 1302
rect 982 1288 986 1292
rect 1014 1288 1018 1292
rect 1190 1288 1194 1292
rect 1230 1288 1234 1292
rect 1262 1288 1266 1292
rect 1318 1288 1322 1292
rect 1334 1288 1338 1292
rect 502 1278 506 1282
rect 518 1278 522 1282
rect 734 1278 738 1282
rect 750 1278 754 1282
rect 838 1278 842 1282
rect 1302 1278 1306 1282
rect 86 1218 90 1222
rect 230 1258 234 1262
rect 294 1258 298 1262
rect 190 1238 194 1242
rect 85 1158 89 1162
rect 278 1248 282 1252
rect 294 1238 298 1242
rect 254 1218 258 1222
rect 102 1138 106 1142
rect 166 1138 170 1142
rect 6 888 10 892
rect 182 1128 186 1132
rect 86 1078 90 1082
rect 334 1158 338 1162
rect 270 1128 274 1132
rect 222 1088 226 1092
rect 302 1108 306 1112
rect 302 1098 306 1102
rect 326 1148 330 1152
rect 342 1148 346 1152
rect 310 1088 314 1092
rect 470 1258 474 1262
rect 398 1188 402 1192
rect 366 1138 370 1142
rect 442 1203 446 1207
rect 449 1203 453 1207
rect 534 1208 538 1212
rect 470 1188 474 1192
rect 478 1168 482 1172
rect 406 1148 410 1152
rect 422 1148 426 1152
rect 534 1158 538 1162
rect 494 1138 498 1142
rect 358 1128 362 1132
rect 374 1128 378 1132
rect 342 1118 346 1122
rect 334 1098 338 1102
rect 334 1088 338 1092
rect 142 1068 146 1072
rect 214 1068 218 1072
rect 238 1068 242 1072
rect 286 1068 290 1072
rect 294 1068 298 1072
rect 214 1058 218 1062
rect 198 1048 202 1052
rect 270 1058 274 1062
rect 286 1058 290 1062
rect 246 1038 250 1042
rect 342 1068 346 1072
rect 334 1058 338 1062
rect 342 1058 346 1062
rect 366 1118 370 1122
rect 310 1048 314 1052
rect 302 1028 306 1032
rect 382 1068 386 1072
rect 502 1068 506 1072
rect 382 1048 386 1052
rect 414 1058 418 1062
rect 590 1208 594 1212
rect 582 1158 586 1162
rect 606 1128 610 1132
rect 582 1088 586 1092
rect 518 1048 522 1052
rect 390 1038 394 1042
rect 398 1038 402 1042
rect 302 958 306 962
rect 166 948 170 952
rect 190 948 194 952
rect 382 948 386 952
rect 110 928 114 932
rect 94 908 98 912
rect 118 908 122 912
rect 102 878 106 882
rect 30 858 34 862
rect 46 858 50 862
rect 102 858 106 862
rect 62 848 66 852
rect 158 868 162 872
rect 118 848 122 852
rect 110 808 114 812
rect 222 878 226 882
rect 230 878 234 882
rect 318 928 322 932
rect 342 928 346 932
rect 358 928 362 932
rect 374 928 378 932
rect 302 918 306 922
rect 262 908 266 912
rect 286 908 290 912
rect 262 878 266 882
rect 14 768 18 772
rect 110 768 114 772
rect 198 768 202 772
rect 6 718 10 722
rect 86 758 90 762
rect 246 798 250 802
rect 126 758 130 762
rect 150 758 154 762
rect 222 758 226 762
rect 238 758 242 762
rect 126 748 130 752
rect 14 708 18 712
rect 6 488 10 492
rect 134 688 138 692
rect 158 688 162 692
rect 70 678 74 682
rect 86 678 90 682
rect 70 548 74 552
rect 278 868 282 872
rect 334 918 338 922
rect 334 898 338 902
rect 294 858 298 862
rect 430 1028 434 1032
rect 414 948 418 952
rect 422 948 426 952
rect 478 1008 482 1012
rect 442 1003 446 1007
rect 449 1003 453 1007
rect 438 978 442 982
rect 534 968 538 972
rect 478 948 482 952
rect 494 948 498 952
rect 526 948 530 952
rect 518 938 522 942
rect 342 868 346 872
rect 358 838 362 842
rect 310 808 314 812
rect 286 798 290 802
rect 270 768 274 772
rect 406 798 410 802
rect 398 788 402 792
rect 406 788 410 792
rect 470 918 474 922
rect 494 918 498 922
rect 430 898 434 902
rect 422 778 426 782
rect 390 758 394 762
rect 246 748 250 752
rect 262 748 266 752
rect 334 748 338 752
rect 390 748 394 752
rect 230 738 234 742
rect 486 888 490 892
rect 574 1048 578 1052
rect 686 1258 690 1262
rect 702 1258 706 1262
rect 718 1258 722 1262
rect 734 1188 738 1192
rect 718 1158 722 1162
rect 726 1158 730 1162
rect 622 1138 626 1142
rect 670 1148 674 1152
rect 678 1138 682 1142
rect 742 1178 746 1182
rect 782 1168 786 1172
rect 790 1158 794 1162
rect 710 1148 714 1152
rect 758 1148 762 1152
rect 774 1148 778 1152
rect 798 1148 802 1152
rect 694 1128 698 1132
rect 694 1108 698 1112
rect 646 1088 650 1092
rect 670 1088 674 1092
rect 614 1068 618 1072
rect 590 1058 594 1062
rect 614 1058 618 1062
rect 694 1078 698 1082
rect 734 1138 738 1142
rect 782 1138 786 1142
rect 822 1138 826 1142
rect 646 1058 650 1062
rect 670 1058 674 1062
rect 702 1058 706 1062
rect 726 1058 730 1062
rect 646 1038 650 1042
rect 702 1028 706 1032
rect 638 1008 642 1012
rect 718 998 722 1002
rect 622 988 626 992
rect 718 988 722 992
rect 758 1128 762 1132
rect 798 1128 802 1132
rect 830 1108 834 1112
rect 1078 1268 1082 1272
rect 910 1248 914 1252
rect 942 1218 946 1222
rect 854 1208 858 1212
rect 870 1208 874 1212
rect 862 1178 866 1182
rect 846 1158 850 1162
rect 854 1158 858 1162
rect 925 1148 929 1152
rect 934 1148 938 1152
rect 846 1138 850 1142
rect 862 1118 866 1122
rect 838 1098 842 1102
rect 750 1078 754 1082
rect 790 1078 794 1082
rect 878 1078 882 1082
rect 742 1058 746 1062
rect 766 1058 770 1062
rect 774 1038 778 1042
rect 734 1028 738 1032
rect 862 1068 866 1072
rect 862 1058 866 1062
rect 822 1048 826 1052
rect 830 1008 834 1012
rect 910 1008 914 1012
rect 838 988 842 992
rect 566 978 570 982
rect 566 958 570 962
rect 710 968 714 972
rect 1038 1248 1042 1252
rect 1006 1218 1010 1222
rect 1070 1218 1074 1222
rect 1254 1268 1258 1272
rect 958 1148 962 1152
rect 1022 1128 1026 1132
rect 1006 1118 1010 1122
rect 1006 1108 1010 1112
rect 1030 1108 1034 1112
rect 962 1103 966 1107
rect 969 1103 973 1107
rect 1062 1098 1066 1102
rect 950 1088 954 1092
rect 966 1088 970 1092
rect 1054 1078 1058 1082
rect 950 1068 954 1072
rect 1006 1058 1010 1062
rect 958 1048 962 1052
rect 918 988 922 992
rect 910 968 914 972
rect 822 958 826 962
rect 846 958 850 962
rect 886 958 890 962
rect 726 948 730 952
rect 742 948 746 952
rect 782 948 786 952
rect 798 948 802 952
rect 606 928 610 932
rect 742 928 746 932
rect 622 908 626 912
rect 654 908 658 912
rect 766 938 770 942
rect 758 928 762 932
rect 750 898 754 902
rect 718 888 722 892
rect 742 888 746 892
rect 598 878 602 882
rect 558 868 562 872
rect 502 858 506 862
rect 550 858 554 862
rect 478 818 482 822
rect 442 803 446 807
rect 449 803 453 807
rect 582 858 586 862
rect 526 788 530 792
rect 438 768 442 772
rect 438 758 442 762
rect 462 758 466 762
rect 318 728 322 732
rect 422 698 426 702
rect 486 698 490 702
rect 574 758 578 762
rect 518 708 522 712
rect 518 698 522 702
rect 198 688 202 692
rect 222 688 226 692
rect 246 688 250 692
rect 342 688 346 692
rect 502 688 506 692
rect 182 638 186 642
rect 174 588 178 592
rect 222 668 226 672
rect 390 678 394 682
rect 454 678 458 682
rect 534 678 538 682
rect 566 678 570 682
rect 222 638 226 642
rect 254 638 258 642
rect 214 618 218 622
rect 190 588 194 592
rect 326 648 330 652
rect 502 668 506 672
rect 510 668 514 672
rect 574 668 578 672
rect 590 718 594 722
rect 638 808 642 812
rect 678 808 682 812
rect 710 768 714 772
rect 670 758 674 762
rect 606 748 610 752
rect 710 748 714 752
rect 598 678 602 682
rect 694 738 698 742
rect 782 898 786 902
rect 814 928 818 932
rect 806 898 810 902
rect 790 878 794 882
rect 798 868 802 872
rect 734 848 738 852
rect 742 838 746 842
rect 758 848 762 852
rect 814 848 818 852
rect 854 948 858 952
rect 774 838 778 842
rect 822 838 826 842
rect 862 918 866 922
rect 966 1018 970 1022
rect 950 958 954 962
rect 1134 1208 1138 1212
rect 1190 1208 1194 1212
rect 1126 1138 1130 1142
rect 1086 1108 1090 1112
rect 1070 1078 1074 1082
rect 1118 1098 1122 1102
rect 1142 1098 1146 1102
rect 1158 1088 1162 1092
rect 1078 1058 1082 1062
rect 1118 1068 1122 1072
rect 1150 1068 1154 1072
rect 1102 1048 1106 1052
rect 1086 1028 1090 1032
rect 1094 1028 1098 1032
rect 1022 1018 1026 1022
rect 1062 1018 1066 1022
rect 990 1008 994 1012
rect 1030 1008 1034 1012
rect 990 988 994 992
rect 1038 998 1042 1002
rect 1086 978 1090 982
rect 1054 968 1058 972
rect 1118 1048 1122 1052
rect 1110 1008 1114 1012
rect 1398 1298 1402 1302
rect 1414 1298 1418 1302
rect 1430 1298 1434 1302
rect 1382 1288 1386 1292
rect 1422 1278 1426 1282
rect 1350 1228 1354 1232
rect 1358 1168 1362 1172
rect 1270 1128 1274 1132
rect 1286 1088 1290 1092
rect 1302 1088 1306 1092
rect 1230 1078 1234 1082
rect 1398 1178 1402 1182
rect 1406 1128 1410 1132
rect 1438 1238 1442 1242
rect 1406 1118 1410 1122
rect 1422 1118 1426 1122
rect 1382 1098 1386 1102
rect 1158 1058 1162 1062
rect 1230 1058 1234 1062
rect 1342 1058 1346 1062
rect 1438 1058 1442 1062
rect 1134 988 1138 992
rect 1382 1028 1386 1032
rect 1326 1008 1330 1012
rect 1438 1038 1442 1042
rect 1438 1008 1442 1012
rect 1390 988 1394 992
rect 1398 988 1402 992
rect 1190 978 1194 982
rect 1262 978 1266 982
rect 1094 968 1098 972
rect 950 948 954 952
rect 1006 948 1010 952
rect 1046 948 1050 952
rect 950 938 954 942
rect 958 928 962 932
rect 966 918 970 922
rect 910 908 914 912
rect 962 903 966 907
rect 969 903 973 907
rect 886 898 890 902
rect 910 888 914 892
rect 982 878 986 882
rect 846 858 850 862
rect 862 858 866 862
rect 862 848 866 852
rect 870 838 874 842
rect 742 778 746 782
rect 750 778 754 782
rect 734 758 738 762
rect 774 768 778 772
rect 830 768 834 772
rect 854 768 858 772
rect 870 768 874 772
rect 830 758 834 762
rect 774 738 778 742
rect 798 748 802 752
rect 750 718 754 722
rect 782 718 786 722
rect 686 688 690 692
rect 726 688 730 692
rect 742 678 746 682
rect 518 658 522 662
rect 550 658 554 662
rect 582 658 586 662
rect 510 638 514 642
rect 438 628 442 632
rect 442 603 446 607
rect 449 603 453 607
rect 174 538 178 542
rect 590 598 594 602
rect 726 638 730 642
rect 614 608 618 612
rect 638 588 642 592
rect 702 608 706 612
rect 630 578 634 582
rect 646 578 650 582
rect 686 578 690 582
rect 502 558 506 562
rect 606 558 610 562
rect 542 548 546 552
rect 486 538 490 542
rect 230 528 234 532
rect 246 528 250 532
rect 294 528 298 532
rect 310 528 314 532
rect 86 518 90 522
rect 118 508 122 512
rect 102 478 106 482
rect 294 508 298 512
rect 310 508 314 512
rect 22 458 26 462
rect 46 458 50 462
rect 158 458 162 462
rect 222 458 226 462
rect 278 458 282 462
rect 206 428 210 432
rect 206 358 210 362
rect 22 348 26 352
rect 46 348 50 352
rect 198 348 202 352
rect 222 348 226 352
rect 278 348 282 352
rect 102 328 106 332
rect 86 308 90 312
rect 118 308 122 312
rect 70 258 74 262
rect 62 218 66 222
rect 14 138 18 142
rect 30 138 34 142
rect 558 518 562 522
rect 446 508 450 512
rect 478 498 482 502
rect 590 498 594 502
rect 598 498 602 502
rect 422 478 426 482
rect 414 458 418 462
rect 382 448 386 452
rect 374 438 378 442
rect 390 428 394 432
rect 422 418 426 422
rect 398 358 402 362
rect 334 348 338 352
rect 262 308 266 312
rect 294 308 298 312
rect 246 278 250 282
rect 126 258 130 262
rect 190 258 194 262
rect 174 238 178 242
rect 302 248 306 252
rect 262 218 266 222
rect 238 158 242 162
rect 142 148 146 152
rect 294 148 298 152
rect 86 128 90 132
rect 158 118 162 122
rect 318 188 322 192
rect 310 158 314 162
rect 422 348 426 352
rect 526 488 530 492
rect 558 478 562 482
rect 614 478 618 482
rect 494 468 498 472
rect 470 458 474 462
rect 486 458 490 462
rect 442 403 446 407
rect 449 403 453 407
rect 478 418 482 422
rect 470 368 474 372
rect 446 338 450 342
rect 454 338 458 342
rect 390 298 394 302
rect 406 288 410 292
rect 398 278 402 282
rect 422 268 426 272
rect 374 258 378 262
rect 414 258 418 262
rect 438 308 442 312
rect 662 568 666 572
rect 694 568 698 572
rect 782 628 786 632
rect 806 738 810 742
rect 798 728 802 732
rect 814 698 818 702
rect 942 868 946 872
rect 902 858 906 862
rect 918 858 922 862
rect 886 768 890 772
rect 862 758 866 762
rect 878 738 882 742
rect 870 718 874 722
rect 854 698 858 702
rect 798 678 802 682
rect 830 678 834 682
rect 798 658 802 662
rect 830 658 834 662
rect 790 578 794 582
rect 734 568 738 572
rect 822 648 826 652
rect 830 618 834 622
rect 854 668 858 672
rect 910 738 914 742
rect 894 708 898 712
rect 910 708 914 712
rect 934 768 938 772
rect 974 858 978 862
rect 966 818 970 822
rect 966 758 970 762
rect 942 748 946 752
rect 950 728 954 732
rect 886 698 890 702
rect 962 703 966 707
rect 969 703 973 707
rect 1438 968 1442 972
rect 1310 948 1314 952
rect 1150 938 1154 942
rect 1190 938 1194 942
rect 1134 928 1138 932
rect 1062 918 1066 922
rect 1134 918 1138 922
rect 1022 908 1026 912
rect 1070 908 1074 912
rect 1014 888 1018 892
rect 1006 878 1010 882
rect 1046 878 1050 882
rect 1022 868 1026 872
rect 1046 868 1050 872
rect 1054 858 1058 862
rect 1006 848 1010 852
rect 998 768 1002 772
rect 990 738 994 742
rect 982 698 986 702
rect 1126 888 1130 892
rect 1158 878 1162 882
rect 1174 878 1178 882
rect 1086 858 1090 862
rect 1102 858 1106 862
rect 1118 848 1122 852
rect 1070 778 1074 782
rect 1222 918 1226 922
rect 1230 888 1234 892
rect 1198 868 1202 872
rect 1246 868 1250 872
rect 1326 928 1330 932
rect 1166 858 1170 862
rect 1110 838 1114 842
rect 1126 838 1130 842
rect 1126 828 1130 832
rect 1142 828 1146 832
rect 1174 828 1178 832
rect 1054 748 1058 752
rect 1006 718 1010 722
rect 1046 718 1050 722
rect 1142 818 1146 822
rect 1190 838 1194 842
rect 1182 818 1186 822
rect 1182 808 1186 812
rect 1150 768 1154 772
rect 1094 758 1098 762
rect 1086 748 1090 752
rect 1110 738 1114 742
rect 1102 728 1106 732
rect 1142 738 1146 742
rect 1166 738 1170 742
rect 1134 718 1138 722
rect 926 688 930 692
rect 998 688 1002 692
rect 1030 688 1034 692
rect 1118 688 1122 692
rect 918 678 922 682
rect 950 678 954 682
rect 1014 678 1018 682
rect 1038 678 1042 682
rect 878 668 882 672
rect 894 668 898 672
rect 934 668 938 672
rect 902 658 906 662
rect 854 648 858 652
rect 862 628 866 632
rect 846 558 850 562
rect 774 548 778 552
rect 782 548 786 552
rect 662 498 666 502
rect 702 538 706 542
rect 790 538 794 542
rect 798 538 802 542
rect 686 528 690 532
rect 750 528 754 532
rect 670 488 674 492
rect 678 488 682 492
rect 646 478 650 482
rect 678 478 682 482
rect 526 458 530 462
rect 582 458 586 462
rect 598 458 602 462
rect 630 458 634 462
rect 518 448 522 452
rect 566 448 570 452
rect 502 408 506 412
rect 518 398 522 402
rect 526 388 530 392
rect 486 358 490 362
rect 470 278 474 282
rect 510 348 514 352
rect 526 338 530 342
rect 582 418 586 422
rect 566 388 570 392
rect 630 438 634 442
rect 670 468 674 472
rect 678 458 682 462
rect 654 438 658 442
rect 622 428 626 432
rect 654 418 658 422
rect 606 398 610 402
rect 654 398 658 402
rect 566 358 570 362
rect 574 358 578 362
rect 494 328 498 332
rect 518 328 522 332
rect 534 328 538 332
rect 494 308 498 312
rect 614 358 618 362
rect 550 348 554 352
rect 566 348 570 352
rect 678 348 682 352
rect 630 338 634 342
rect 630 328 634 332
rect 558 318 562 322
rect 590 318 594 322
rect 622 318 626 322
rect 526 298 530 302
rect 542 298 546 302
rect 494 278 498 282
rect 502 278 506 282
rect 478 268 482 272
rect 454 248 458 252
rect 478 248 482 252
rect 342 218 346 222
rect 442 203 446 207
rect 449 203 453 207
rect 350 188 354 192
rect 374 188 378 192
rect 446 188 450 192
rect 366 178 370 182
rect 398 178 402 182
rect 438 168 442 172
rect 422 158 426 162
rect 374 148 378 152
rect 390 148 394 152
rect 510 268 514 272
rect 542 268 546 272
rect 598 288 602 292
rect 614 288 618 292
rect 582 268 586 272
rect 606 268 610 272
rect 542 238 546 242
rect 542 228 546 232
rect 534 198 538 202
rect 510 178 514 182
rect 510 168 514 172
rect 462 148 466 152
rect 478 148 482 152
rect 406 138 410 142
rect 486 138 490 142
rect 414 128 418 132
rect 430 128 434 132
rect 374 118 378 122
rect 158 98 162 102
rect 182 98 186 102
rect 198 98 202 102
rect 222 98 226 102
rect 326 98 330 102
rect 166 78 170 82
rect 318 88 322 92
rect 286 78 290 82
rect 294 68 298 72
rect 398 88 402 92
rect 422 88 426 92
rect 350 78 354 82
rect 454 78 458 82
rect 358 68 362 72
rect 430 68 434 72
rect 478 128 482 132
rect 494 118 498 122
rect 502 98 506 102
rect 486 88 490 92
rect 478 78 482 82
rect 486 68 490 72
rect 302 58 306 62
rect 366 58 370 62
rect 390 58 394 62
rect 406 58 410 62
rect 470 58 474 62
rect 574 238 578 242
rect 590 238 594 242
rect 566 228 570 232
rect 582 228 586 232
rect 558 218 562 222
rect 558 178 562 182
rect 550 138 554 142
rect 630 298 634 302
rect 750 518 754 522
rect 774 528 778 532
rect 774 508 778 512
rect 774 498 778 502
rect 774 488 778 492
rect 758 478 762 482
rect 790 478 794 482
rect 798 478 802 482
rect 1006 668 1010 672
rect 990 658 994 662
rect 1198 828 1202 832
rect 1230 838 1234 842
rect 1238 828 1242 832
rect 1310 848 1314 852
rect 1214 808 1218 812
rect 1398 858 1402 862
rect 1422 858 1426 862
rect 1326 808 1330 812
rect 1342 808 1346 812
rect 1206 748 1210 752
rect 1198 718 1202 722
rect 1206 718 1210 722
rect 1174 708 1178 712
rect 1190 708 1194 712
rect 1174 698 1178 702
rect 1046 658 1050 662
rect 1078 658 1082 662
rect 934 648 938 652
rect 1062 648 1066 652
rect 1094 648 1098 652
rect 926 618 930 622
rect 1158 618 1162 622
rect 918 598 922 602
rect 998 598 1002 602
rect 902 548 906 552
rect 1070 588 1074 592
rect 1006 538 1010 542
rect 870 528 874 532
rect 1038 528 1042 532
rect 830 508 834 512
rect 962 503 966 507
rect 969 503 973 507
rect 838 498 842 502
rect 902 498 906 502
rect 926 498 930 502
rect 726 468 730 472
rect 734 468 738 472
rect 750 468 754 472
rect 774 468 778 472
rect 814 468 818 472
rect 694 458 698 462
rect 702 448 706 452
rect 694 428 698 432
rect 694 398 698 402
rect 878 488 882 492
rect 918 478 922 482
rect 886 468 890 472
rect 966 488 970 492
rect 1022 488 1026 492
rect 1046 488 1050 492
rect 934 478 938 482
rect 822 458 826 462
rect 830 458 834 462
rect 878 458 882 462
rect 894 458 898 462
rect 910 458 914 462
rect 742 448 746 452
rect 766 448 770 452
rect 734 428 738 432
rect 758 428 762 432
rect 734 408 738 412
rect 726 398 730 402
rect 710 388 714 392
rect 702 378 706 382
rect 774 388 778 392
rect 758 368 762 372
rect 742 358 746 362
rect 710 348 714 352
rect 766 358 770 362
rect 790 368 794 372
rect 814 398 818 402
rect 790 358 794 362
rect 806 358 810 362
rect 782 348 786 352
rect 702 328 706 332
rect 646 278 650 282
rect 630 248 634 252
rect 630 228 634 232
rect 678 288 682 292
rect 662 258 666 262
rect 646 248 650 252
rect 638 198 642 202
rect 662 198 666 202
rect 694 308 698 312
rect 726 298 730 302
rect 750 298 754 302
rect 774 318 778 322
rect 790 338 794 342
rect 782 308 786 312
rect 758 278 762 282
rect 718 268 722 272
rect 734 248 738 252
rect 702 238 706 242
rect 686 218 690 222
rect 686 178 690 182
rect 726 218 730 222
rect 734 188 738 192
rect 606 148 610 152
rect 638 148 642 152
rect 654 148 658 152
rect 670 148 674 152
rect 718 148 722 152
rect 590 138 594 142
rect 614 118 618 122
rect 582 98 586 102
rect 558 88 562 92
rect 518 78 522 82
rect 542 78 546 82
rect 518 68 522 72
rect 406 48 410 52
rect 494 48 498 52
rect 622 88 626 92
rect 646 88 650 92
rect 590 78 594 82
rect 574 68 578 72
rect 558 58 562 62
rect 606 58 610 62
rect 638 58 642 62
rect 694 138 698 142
rect 734 148 738 152
rect 862 448 866 452
rect 926 448 930 452
rect 886 398 890 402
rect 822 358 826 362
rect 846 358 850 362
rect 870 358 874 362
rect 918 368 922 372
rect 902 358 906 362
rect 822 338 826 342
rect 878 338 882 342
rect 822 328 826 332
rect 806 318 810 322
rect 830 318 834 322
rect 798 308 802 312
rect 806 298 810 302
rect 822 298 826 302
rect 838 308 842 312
rect 862 298 866 302
rect 886 298 890 302
rect 862 268 866 272
rect 878 268 882 272
rect 798 228 802 232
rect 798 198 802 202
rect 822 248 826 252
rect 838 248 842 252
rect 830 238 834 242
rect 846 218 850 222
rect 854 198 858 202
rect 878 228 882 232
rect 862 148 866 152
rect 862 138 866 142
rect 910 338 914 342
rect 902 328 906 332
rect 958 468 962 472
rect 1006 468 1010 472
rect 1030 478 1034 482
rect 982 458 986 462
rect 998 458 1002 462
rect 974 388 978 392
rect 966 368 970 372
rect 934 308 938 312
rect 942 298 946 302
rect 934 278 938 282
rect 902 268 906 272
rect 910 228 914 232
rect 902 218 906 222
rect 894 208 898 212
rect 962 303 966 307
rect 969 303 973 307
rect 1078 578 1082 582
rect 1062 548 1066 552
rect 1054 468 1058 472
rect 1110 568 1114 572
rect 1182 688 1186 692
rect 1182 668 1186 672
rect 1238 618 1242 622
rect 1326 708 1330 712
rect 1342 708 1346 712
rect 1358 708 1362 712
rect 1382 708 1386 712
rect 1286 628 1290 632
rect 1238 598 1242 602
rect 1262 598 1266 602
rect 1110 548 1114 552
rect 1150 548 1154 552
rect 1238 548 1242 552
rect 1094 518 1098 522
rect 1110 518 1114 522
rect 1086 478 1090 482
rect 1094 478 1098 482
rect 1054 438 1058 442
rect 1070 438 1074 442
rect 1134 538 1138 542
rect 1150 528 1154 532
rect 1126 488 1130 492
rect 1190 538 1194 542
rect 1158 518 1162 522
rect 1190 498 1194 502
rect 1214 488 1218 492
rect 1142 478 1146 482
rect 1150 478 1154 482
rect 1166 478 1170 482
rect 1198 478 1202 482
rect 1278 538 1282 542
rect 1326 528 1330 532
rect 1326 518 1330 522
rect 1294 488 1298 492
rect 1254 478 1258 482
rect 1262 478 1266 482
rect 1270 478 1274 482
rect 1366 528 1370 532
rect 1438 648 1442 652
rect 1414 558 1418 562
rect 1406 478 1410 482
rect 1142 468 1146 472
rect 1158 468 1162 472
rect 1182 468 1186 472
rect 1254 468 1258 472
rect 1350 468 1354 472
rect 1166 458 1170 462
rect 1222 458 1226 462
rect 1230 458 1234 462
rect 1238 458 1242 462
rect 1262 458 1266 462
rect 1190 448 1194 452
rect 1102 438 1106 442
rect 1126 438 1130 442
rect 1078 428 1082 432
rect 1086 428 1090 432
rect 1014 378 1018 382
rect 1014 358 1018 362
rect 982 288 986 292
rect 974 278 978 282
rect 1062 358 1066 362
rect 1022 338 1026 342
rect 1046 338 1050 342
rect 1086 358 1090 362
rect 1118 388 1122 392
rect 1102 348 1106 352
rect 1142 368 1146 372
rect 1150 358 1154 362
rect 1182 358 1186 362
rect 1190 358 1194 362
rect 1214 448 1218 452
rect 1358 448 1362 452
rect 1302 438 1306 442
rect 1230 368 1234 372
rect 1414 448 1418 452
rect 1406 358 1410 362
rect 1206 348 1210 352
rect 1238 348 1242 352
rect 1270 348 1274 352
rect 1398 348 1402 352
rect 1070 338 1074 342
rect 1102 338 1106 342
rect 1198 338 1202 342
rect 1222 338 1226 342
rect 1062 328 1066 332
rect 1038 318 1042 322
rect 1102 318 1106 322
rect 1038 308 1042 312
rect 942 258 946 262
rect 990 258 994 262
rect 926 198 930 202
rect 958 198 962 202
rect 926 178 930 182
rect 910 158 914 162
rect 966 168 970 172
rect 934 158 938 162
rect 958 158 962 162
rect 918 148 922 152
rect 926 148 930 152
rect 950 148 954 152
rect 894 138 898 142
rect 926 138 930 142
rect 910 128 914 132
rect 934 128 938 132
rect 854 98 858 102
rect 814 88 818 92
rect 702 78 706 82
rect 926 78 930 82
rect 966 138 970 142
rect 962 103 966 107
rect 969 103 973 107
rect 958 78 962 82
rect 694 68 698 72
rect 734 68 738 72
rect 878 68 882 72
rect 718 58 722 62
rect 686 48 690 52
rect 534 38 538 42
rect 646 38 650 42
rect 910 58 914 62
rect 1006 218 1010 222
rect 1030 218 1034 222
rect 1022 208 1026 212
rect 1014 198 1018 202
rect 1014 138 1018 142
rect 1014 128 1018 132
rect 990 68 994 72
rect 950 58 954 62
rect 1030 148 1034 152
rect 1030 118 1034 122
rect 1134 328 1138 332
rect 1174 328 1178 332
rect 1118 278 1122 282
rect 1102 268 1106 272
rect 1174 268 1178 272
rect 1054 258 1058 262
rect 1046 248 1050 252
rect 1118 258 1122 262
rect 1182 258 1186 262
rect 1102 238 1106 242
rect 1054 228 1058 232
rect 1062 148 1066 152
rect 1054 138 1058 142
rect 1046 128 1050 132
rect 1134 198 1138 202
rect 1118 178 1122 182
rect 1406 338 1410 342
rect 1334 328 1338 332
rect 1278 318 1282 322
rect 1318 318 1322 322
rect 1374 318 1378 322
rect 1238 268 1242 272
rect 1294 258 1298 262
rect 1238 198 1242 202
rect 1302 198 1306 202
rect 1342 198 1346 202
rect 1374 198 1378 202
rect 1150 178 1154 182
rect 1198 178 1202 182
rect 1214 178 1218 182
rect 1230 178 1234 182
rect 1238 178 1242 182
rect 1126 158 1130 162
rect 1198 168 1202 172
rect 1182 158 1186 162
rect 1214 168 1218 172
rect 1254 148 1258 152
rect 1134 138 1138 142
rect 1214 138 1218 142
rect 1078 128 1082 132
rect 1110 128 1114 132
rect 1078 98 1082 102
rect 1086 88 1090 92
rect 1118 78 1122 82
rect 1086 68 1090 72
rect 1110 68 1114 72
rect 1126 68 1130 72
rect 1102 58 1106 62
rect 1142 128 1146 132
rect 1254 118 1258 122
rect 1238 108 1242 112
rect 1142 98 1146 102
rect 1358 148 1362 152
rect 1342 108 1346 112
rect 1366 108 1370 112
rect 1326 98 1330 102
rect 1430 608 1434 612
rect 1438 448 1442 452
rect 1438 348 1442 352
rect 1422 118 1426 122
rect 1438 118 1442 122
rect 1334 88 1338 92
rect 1254 58 1258 62
rect 942 48 946 52
rect 974 48 978 52
rect 982 48 986 52
rect 1094 38 1098 42
rect 1358 48 1362 52
rect 1310 8 1314 12
rect 1334 8 1338 12
rect 1406 8 1410 12
rect 1422 8 1426 12
rect 442 3 446 7
rect 449 3 453 7
<< metal3 >>
rect 1470 1318 1474 1322
rect -26 1308 -22 1312
rect 1470 1311 1473 1318
rect 1462 1308 1473 1311
rect -26 1301 -23 1308
rect 960 1303 962 1307
rect 966 1303 969 1307
rect 974 1303 976 1307
rect -26 1298 30 1301
rect 1002 1298 1006 1301
rect 1210 1298 1270 1301
rect 1282 1298 1286 1301
rect 1306 1298 1350 1301
rect 1362 1298 1366 1301
rect 1378 1298 1382 1301
rect 1394 1298 1398 1301
rect 1410 1298 1414 1301
rect 1426 1298 1430 1301
rect 1462 1301 1465 1308
rect 1442 1298 1465 1301
rect 1470 1298 1474 1302
rect -26 1291 -22 1292
rect -26 1288 38 1291
rect 986 1288 1014 1291
rect 1182 1288 1190 1291
rect 1194 1288 1214 1291
rect 1254 1288 1262 1291
rect 1302 1288 1318 1291
rect 1330 1288 1334 1291
rect 1346 1288 1382 1291
rect 1470 1291 1473 1298
rect 1426 1288 1473 1291
rect 522 1278 734 1281
rect 738 1278 750 1281
rect 1230 1281 1233 1288
rect 1302 1282 1305 1288
rect 842 1278 1081 1281
rect 1230 1278 1262 1281
rect 1470 1281 1474 1282
rect 1426 1278 1474 1281
rect -26 1271 -22 1272
rect 502 1271 505 1278
rect -26 1268 505 1271
rect 1078 1272 1081 1278
rect 1082 1268 1254 1271
rect 234 1258 294 1261
rect 474 1258 478 1261
rect 690 1258 702 1261
rect 714 1258 718 1261
rect 1470 1261 1474 1262
rect 1434 1258 1474 1261
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 282 1248 286 1251
rect 914 1248 1038 1251
rect 194 1238 294 1241
rect 1470 1241 1474 1242
rect 1442 1238 1474 1241
rect 10 1218 14 1221
rect 50 1218 86 1221
rect 90 1218 254 1221
rect 946 1218 1006 1221
rect 1010 1218 1070 1221
rect 1350 1221 1353 1228
rect 1470 1221 1474 1222
rect 1350 1218 1474 1221
rect 538 1208 590 1211
rect 858 1208 870 1211
rect 1138 1208 1190 1211
rect 440 1203 442 1207
rect 446 1203 449 1207
rect 454 1203 456 1207
rect 1470 1201 1474 1202
rect 1410 1198 1474 1201
rect 402 1188 470 1191
rect 474 1188 734 1191
rect 746 1178 750 1181
rect 754 1178 862 1181
rect 1470 1181 1474 1182
rect 1402 1178 1474 1181
rect 482 1168 721 1171
rect 718 1162 721 1168
rect 1362 1168 1422 1171
rect 26 1158 85 1161
rect 338 1158 534 1161
rect 782 1161 785 1168
rect 730 1158 785 1161
rect 794 1158 846 1161
rect 1470 1161 1474 1162
rect 1426 1158 1474 1161
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 18 1148 57 1151
rect 330 1148 342 1151
rect 410 1148 422 1151
rect 582 1151 585 1158
rect 582 1148 670 1151
rect 714 1148 758 1151
rect 766 1148 774 1151
rect 778 1148 798 1151
rect 854 1151 857 1158
rect 854 1148 862 1151
rect 938 1148 958 1151
rect 54 1142 57 1148
rect 106 1138 166 1141
rect 170 1138 366 1141
rect 370 1138 494 1141
rect 626 1138 678 1141
rect 682 1138 734 1141
rect 738 1138 782 1141
rect 926 1141 929 1148
rect 850 1138 929 1141
rect 1470 1141 1474 1142
rect 1130 1138 1273 1141
rect 186 1128 270 1131
rect 274 1128 358 1131
rect 362 1128 374 1131
rect 378 1128 606 1131
rect 610 1128 694 1131
rect 762 1128 798 1131
rect 822 1131 825 1138
rect 1270 1132 1273 1138
rect 1406 1138 1474 1141
rect 1406 1132 1409 1138
rect 822 1128 1022 1131
rect 346 1118 366 1121
rect 866 1118 1006 1121
rect 1410 1118 1422 1121
rect 1470 1121 1474 1122
rect 1442 1118 1474 1121
rect 306 1108 574 1111
rect 698 1108 830 1111
rect 834 1108 886 1111
rect 1002 1108 1006 1111
rect 1034 1108 1086 1111
rect 960 1103 962 1107
rect 966 1103 969 1107
rect 974 1103 976 1107
rect 306 1098 334 1101
rect 834 1098 838 1101
rect 1066 1098 1118 1101
rect 1122 1098 1142 1101
rect 1470 1101 1474 1102
rect 1386 1098 1474 1101
rect 314 1088 334 1091
rect 338 1088 582 1091
rect 586 1088 646 1091
rect 650 1088 670 1091
rect 954 1088 966 1091
rect 970 1088 1158 1091
rect 1290 1088 1302 1091
rect 222 1081 225 1088
rect 90 1078 225 1081
rect 686 1078 694 1081
rect 698 1078 742 1081
rect 754 1078 790 1081
rect 1058 1078 1070 1081
rect 1470 1081 1474 1082
rect 1418 1078 1474 1081
rect 878 1072 881 1078
rect 146 1068 214 1071
rect 242 1068 286 1071
rect 298 1068 342 1071
rect 374 1068 382 1071
rect 386 1068 494 1071
rect 506 1068 614 1071
rect 618 1068 862 1071
rect 866 1068 870 1071
rect 954 1068 1081 1071
rect 1078 1062 1081 1068
rect 1230 1071 1233 1078
rect 1154 1068 1233 1071
rect 218 1058 270 1061
rect 278 1058 286 1061
rect 290 1058 334 1061
rect 346 1058 414 1061
rect 422 1058 590 1061
rect 618 1058 646 1061
rect 674 1058 702 1061
rect 730 1058 742 1061
rect 770 1058 862 1061
rect 962 1058 1006 1061
rect 1118 1061 1121 1068
rect 1118 1058 1158 1061
rect 1234 1058 1342 1061
rect 1470 1061 1474 1062
rect 1442 1058 1474 1061
rect 202 1048 310 1051
rect 422 1051 425 1058
rect 1102 1052 1105 1058
rect 386 1048 425 1051
rect 498 1048 518 1051
rect 578 1048 822 1051
rect 882 1048 958 1051
rect 1122 1048 1126 1051
rect 250 1038 390 1041
rect 402 1038 478 1041
rect 650 1038 774 1041
rect 1470 1041 1474 1042
rect 1442 1038 1474 1041
rect 306 1028 430 1031
rect 434 1028 694 1031
rect 698 1028 702 1031
rect 706 1028 734 1031
rect 746 1028 1086 1031
rect 1098 1028 1166 1031
rect 630 1018 958 1021
rect 970 1018 1022 1021
rect 1026 1018 1062 1021
rect 1382 1021 1385 1028
rect 1470 1021 1474 1022
rect 1382 1018 1474 1021
rect 630 1011 633 1018
rect 482 1008 633 1011
rect 642 1008 830 1011
rect 914 1008 990 1011
rect 1034 1008 1110 1011
rect 1114 1008 1326 1011
rect 1434 1008 1438 1011
rect 440 1003 442 1007
rect 446 1003 449 1007
rect 454 1003 456 1007
rect 722 998 1038 1001
rect 438 988 606 991
rect 610 988 622 991
rect 626 988 718 991
rect 842 988 878 991
rect 922 988 990 991
rect 994 988 1134 991
rect 1170 988 1390 991
rect 1394 988 1398 991
rect 438 982 441 988
rect 570 978 1086 981
rect 1090 978 1190 981
rect 1194 978 1262 981
rect 1438 972 1441 978
rect 538 968 710 971
rect 714 968 910 971
rect 1058 968 1094 971
rect 306 958 566 961
rect 578 958 729 961
rect 826 958 846 961
rect 890 958 950 961
rect 726 952 729 958
rect 170 948 190 951
rect 386 948 414 951
rect 418 948 422 951
rect 482 948 486 951
rect 498 948 526 951
rect 786 948 798 951
rect 954 948 982 951
rect 1010 948 1046 951
rect 742 941 745 948
rect 766 942 769 948
rect 854 942 857 948
rect 522 938 609 941
rect 742 938 750 941
rect 954 938 1137 941
rect 110 932 113 938
rect 606 932 609 938
rect 1134 932 1137 938
rect 1310 941 1313 948
rect 1194 938 1313 941
rect 322 928 342 931
rect 362 928 374 931
rect 746 928 758 931
rect 818 928 958 931
rect 1150 931 1153 938
rect 1150 928 1326 931
rect 282 918 302 921
rect 306 918 334 921
rect 466 918 470 921
rect 498 918 862 921
rect 866 918 966 921
rect 1066 918 1134 921
rect 1226 918 1230 921
rect 98 908 118 911
rect 122 908 262 911
rect 494 911 497 918
rect 290 908 497 911
rect 626 908 654 911
rect 658 908 838 911
rect 850 908 910 911
rect 1026 908 1070 911
rect 960 903 962 907
rect 966 903 969 907
rect 974 903 976 907
rect 338 898 430 901
rect 434 898 750 901
rect 754 898 782 901
rect 810 898 886 901
rect 10 888 14 891
rect 722 888 742 891
rect 746 888 750 891
rect 914 888 1014 891
rect 1118 888 1126 891
rect 1130 888 1230 891
rect 226 878 230 881
rect 486 881 489 888
rect 266 878 598 881
rect 794 878 982 881
rect 1010 878 1046 881
rect 1162 878 1166 881
rect 102 871 105 878
rect 102 868 158 871
rect 502 868 558 871
rect 802 868 862 871
rect 946 868 1022 871
rect 1050 868 1158 871
rect 1174 871 1177 878
rect 1174 868 1198 871
rect 1242 868 1246 871
rect 34 858 46 861
rect 106 858 110 861
rect 278 861 281 868
rect 278 858 294 861
rect 342 861 345 868
rect 298 858 345 861
rect 502 862 505 868
rect 862 862 865 868
rect 554 858 582 861
rect 814 858 846 861
rect 850 858 857 861
rect 906 858 918 861
rect 978 858 1054 861
rect 1090 858 1102 861
rect 1170 858 1334 861
rect 1338 858 1398 861
rect 1402 858 1422 861
rect 814 852 817 858
rect 66 848 118 851
rect 738 848 758 851
rect 858 848 862 851
rect 1010 848 1118 851
rect 1230 848 1310 851
rect 1230 842 1233 848
rect 362 838 742 841
rect 778 838 822 841
rect 874 838 1110 841
rect 1114 838 1126 841
rect 1130 838 1190 841
rect 1106 828 1126 831
rect 1146 828 1174 831
rect 1202 828 1238 831
rect 482 818 486 821
rect 970 818 1126 821
rect 1146 818 1182 821
rect 114 808 310 811
rect 642 808 678 811
rect 1186 808 1214 811
rect 1330 808 1342 811
rect 440 803 442 807
rect 446 803 449 807
rect 454 803 456 807
rect 250 798 286 801
rect 410 798 417 801
rect 402 788 406 791
rect 414 791 417 798
rect 414 788 526 791
rect 530 788 846 791
rect 426 778 441 781
rect 746 778 750 781
rect 754 778 1070 781
rect 438 772 441 778
rect 18 768 110 771
rect 202 768 270 771
rect 778 768 782 771
rect 834 768 854 771
rect 874 768 878 771
rect 890 768 934 771
rect 946 768 998 771
rect 1002 768 1150 771
rect 90 758 126 761
rect 154 758 222 761
rect 242 758 390 761
rect 466 758 526 761
rect 578 758 670 761
rect 710 761 713 768
rect 674 758 713 761
rect 730 758 734 761
rect 786 758 830 761
rect 834 758 862 761
rect 866 758 966 761
rect 130 748 246 751
rect 266 748 334 751
rect 438 751 441 758
rect 394 748 441 751
rect 610 748 614 751
rect 714 748 718 751
rect 802 748 942 751
rect 1058 748 1086 751
rect 1094 751 1097 758
rect 1094 748 1206 751
rect 694 742 697 748
rect 234 738 321 741
rect 778 738 801 741
rect 810 738 878 741
rect 882 738 910 741
rect 994 738 998 741
rect 1002 738 1110 741
rect 1114 738 1142 741
rect 1146 738 1166 741
rect 318 732 321 738
rect 798 732 801 738
rect 806 728 950 731
rect 954 728 1102 731
rect 10 718 590 721
rect 594 718 742 721
rect 754 718 782 721
rect 806 721 809 728
rect 786 718 809 721
rect 866 718 870 721
rect 874 718 1006 721
rect 1010 718 1046 721
rect 1050 718 1134 721
rect 1138 718 1198 721
rect 1202 718 1206 721
rect 18 708 518 711
rect 522 708 710 711
rect 714 708 814 711
rect 898 708 910 711
rect 1178 708 1190 711
rect 1330 708 1342 711
rect 1362 708 1382 711
rect 960 703 962 707
rect 966 703 969 707
rect 974 703 976 707
rect 426 698 486 701
rect 490 698 518 701
rect 530 698 814 701
rect 858 698 886 701
rect 986 698 1174 701
rect 138 688 158 691
rect 162 688 198 691
rect 226 688 246 691
rect 506 688 686 691
rect 930 688 998 691
rect 1002 688 1030 691
rect 1034 688 1118 691
rect 1122 688 1182 691
rect 342 681 345 688
rect 502 682 505 688
rect 90 678 345 681
rect 394 678 454 681
rect 458 678 462 681
rect 538 678 566 681
rect 726 681 729 688
rect 602 678 729 681
rect 802 678 830 681
rect 922 678 934 681
rect 938 678 950 681
rect 954 678 1014 681
rect 1018 678 1038 681
rect 70 671 73 678
rect 70 668 222 671
rect 514 668 574 671
rect 742 671 745 678
rect 894 672 897 678
rect 742 668 798 671
rect 858 668 878 671
rect 938 668 942 671
rect 954 668 1006 671
rect 1010 668 1182 671
rect 502 661 505 668
rect 502 658 518 661
rect 586 658 718 661
rect 802 658 830 661
rect 834 658 902 661
rect 906 658 990 661
rect 994 658 1046 661
rect 1050 658 1078 661
rect 550 651 553 658
rect 330 648 553 651
rect 730 648 822 651
rect 826 648 854 651
rect 858 648 865 651
rect 1066 648 1094 651
rect 1470 651 1474 652
rect 1442 648 1474 651
rect 186 638 222 641
rect 226 638 254 641
rect 258 638 510 641
rect 698 638 726 641
rect 934 641 937 648
rect 730 638 1190 641
rect 786 628 862 631
rect 866 628 1286 631
rect 438 621 441 628
rect 218 618 441 621
rect 466 618 830 621
rect 834 618 926 621
rect 1162 618 1238 621
rect 618 608 702 611
rect 746 608 1430 611
rect 440 603 442 607
rect 446 603 449 607
rect 454 603 456 607
rect 594 598 870 601
rect 874 598 918 601
rect 1242 598 1262 601
rect 998 592 1001 598
rect 178 588 190 591
rect 642 588 857 591
rect 1002 588 1070 591
rect 634 578 646 581
rect 690 578 790 581
rect 854 581 857 588
rect 854 578 1078 581
rect 666 568 694 571
rect 706 568 734 571
rect 738 568 1110 571
rect -26 561 -22 562
rect -26 558 462 561
rect 610 558 774 561
rect 850 558 1414 561
rect 502 552 505 558
rect 774 552 777 558
rect 786 548 801 551
rect 70 541 73 548
rect 70 538 174 541
rect 294 538 486 541
rect 542 541 545 548
rect 798 542 801 548
rect 1066 548 1110 551
rect 1114 548 1150 551
rect 1154 548 1238 551
rect 542 538 702 541
rect 902 541 905 548
rect 902 538 1006 541
rect 1138 538 1190 541
rect 294 532 297 538
rect 790 532 793 538
rect 234 528 246 531
rect 314 528 561 531
rect 690 528 750 531
rect 778 528 782 531
rect 814 528 870 531
rect 1042 528 1118 531
rect 1122 528 1150 531
rect 1278 531 1281 538
rect 1278 528 1326 531
rect 1330 528 1366 531
rect 86 522 89 528
rect 558 522 561 528
rect 814 521 817 528
rect 754 518 817 521
rect 1098 518 1110 521
rect 1114 518 1158 521
rect 1162 518 1326 521
rect 122 508 294 511
rect 298 508 310 511
rect 450 508 774 511
rect 834 508 894 511
rect 960 503 962 507
rect 966 503 969 507
rect 974 503 976 507
rect 482 498 590 501
rect 602 498 662 501
rect 778 498 838 501
rect 906 498 926 501
rect 930 498 934 501
rect 1194 498 1358 501
rect 530 488 670 491
rect 682 488 694 491
rect 698 488 774 491
rect 802 488 878 491
rect 890 488 966 491
rect 1026 488 1046 491
rect 1050 488 1126 491
rect 1218 488 1294 491
rect 6 482 9 488
rect 106 478 422 481
rect 562 478 614 481
rect 618 478 638 481
rect 682 478 758 481
rect 762 478 790 481
rect 802 478 918 481
rect 1034 478 1086 481
rect 1098 478 1142 481
rect 1154 478 1166 481
rect 1202 478 1254 481
rect 1266 478 1270 481
rect 278 468 489 471
rect 278 462 281 468
rect 486 462 489 468
rect 646 471 649 478
rect 646 468 670 471
rect 674 468 726 471
rect 738 468 750 471
rect 778 468 814 471
rect 934 471 937 478
rect 890 468 937 471
rect 962 468 1006 471
rect 1010 468 1054 471
rect 1146 468 1158 471
rect 1186 468 1254 471
rect 1258 468 1350 471
rect 1406 471 1409 478
rect 1354 468 1409 471
rect 26 458 46 461
rect 162 458 222 461
rect 418 458 470 461
rect 494 461 497 468
rect 830 462 833 468
rect 494 458 526 461
rect 586 458 598 461
rect 634 458 678 461
rect 698 458 822 461
rect 834 458 878 461
rect 898 458 902 461
rect 914 458 982 461
rect 1170 458 1222 461
rect 1242 458 1262 461
rect 386 448 518 451
rect 570 448 702 451
rect 746 448 750 451
rect 754 448 766 451
rect 866 448 926 451
rect 998 451 1001 458
rect 998 448 1190 451
rect 1194 448 1214 451
rect 1230 451 1233 458
rect 1230 448 1358 451
rect 1418 448 1422 451
rect 1470 451 1474 452
rect 1442 448 1474 451
rect 378 438 630 441
rect 658 438 790 441
rect 1058 438 1070 441
rect 1074 438 1102 441
rect 1130 438 1302 441
rect 210 428 390 431
rect 394 428 622 431
rect 626 428 694 431
rect 730 428 734 431
rect 762 428 1078 431
rect 1082 428 1086 431
rect 426 418 478 421
rect 482 418 582 421
rect 586 418 654 421
rect 506 408 734 411
rect 440 403 442 407
rect 446 403 449 407
rect 454 403 456 407
rect 522 398 606 401
rect 610 398 654 401
rect 658 398 694 401
rect 730 398 814 401
rect 818 398 886 401
rect 1118 392 1121 398
rect 530 388 566 391
rect 714 388 774 391
rect 818 388 974 391
rect 706 378 1014 381
rect 474 368 758 371
rect 786 368 790 371
rect 794 368 801 371
rect 970 368 1142 371
rect 1146 368 1230 371
rect 918 362 921 368
rect 210 358 398 361
rect 490 358 566 361
rect 578 358 614 361
rect 746 358 766 361
rect 794 358 798 361
rect 802 358 806 361
rect 826 358 846 361
rect 850 358 870 361
rect 906 358 910 361
rect 1018 358 1062 361
rect 1090 358 1150 361
rect 1154 358 1182 361
rect 1194 358 1198 361
rect 1410 358 1422 361
rect 26 348 46 351
rect 202 348 222 351
rect 338 348 422 351
rect 426 348 510 351
rect 554 348 566 351
rect 698 348 710 351
rect 778 348 782 351
rect 786 348 1073 351
rect 1106 348 1206 351
rect 1210 348 1214 351
rect 1242 348 1270 351
rect 1362 348 1390 351
rect 1394 348 1398 351
rect 1470 351 1474 352
rect 1442 348 1474 351
rect 278 342 281 348
rect 450 338 454 341
rect 458 338 526 341
rect 678 341 681 348
rect 1070 342 1073 348
rect 634 338 681 341
rect 722 338 790 341
rect 818 338 822 341
rect 882 338 910 341
rect 1026 338 1046 341
rect 1106 338 1134 341
rect 1138 338 1198 341
rect 1202 338 1222 341
rect 1410 338 1414 341
rect 102 332 105 338
rect 522 328 534 331
rect 546 328 630 331
rect 642 328 702 331
rect 786 328 822 331
rect 906 328 1062 331
rect 1066 328 1134 331
rect 1178 328 1334 331
rect 494 322 497 328
rect 562 318 590 321
rect 626 318 734 321
rect 778 318 806 321
rect 834 318 1038 321
rect 1106 318 1278 321
rect 1282 318 1318 321
rect 1322 318 1374 321
rect 90 308 118 311
rect 266 308 294 311
rect 442 308 494 311
rect 506 308 694 311
rect 698 308 782 311
rect 802 308 838 311
rect 930 308 934 311
rect 1042 308 1230 311
rect 960 303 962 307
rect 966 303 969 307
rect 974 303 976 307
rect 394 298 526 301
rect 530 298 542 301
rect 546 298 630 301
rect 706 298 726 301
rect 754 298 790 301
rect 794 298 806 301
rect 826 298 830 301
rect 850 298 862 301
rect 890 298 942 301
rect 410 288 497 291
rect 602 288 614 291
rect 618 288 678 291
rect 682 288 982 291
rect 494 282 497 288
rect 402 278 470 281
rect 506 278 646 281
rect 650 278 758 281
rect 762 278 822 281
rect 938 278 974 281
rect 1102 278 1118 281
rect 246 271 249 278
rect 1102 272 1105 278
rect 246 268 422 271
rect 482 268 510 271
rect 518 268 542 271
rect 586 268 606 271
rect 626 268 718 271
rect 866 268 873 271
rect 882 268 902 271
rect 1178 268 1238 271
rect 70 262 73 268
rect 130 258 190 261
rect 378 258 414 261
rect 518 261 521 268
rect 1118 262 1121 268
rect 418 258 521 261
rect 538 258 662 261
rect 826 258 942 261
rect 994 258 1054 261
rect 1186 258 1294 261
rect 306 248 454 251
rect 482 248 593 251
rect 634 248 646 251
rect 738 248 822 251
rect 842 248 1046 251
rect 590 242 593 248
rect 178 238 534 241
rect 546 238 574 241
rect 706 238 718 241
rect 722 238 830 241
rect 834 238 1102 241
rect 342 228 542 231
rect 546 228 566 231
rect 570 228 582 231
rect 634 228 750 231
rect 802 228 878 231
rect 882 228 910 231
rect 914 228 1054 231
rect 342 222 345 228
rect 66 218 262 221
rect 562 218 566 221
rect 690 218 726 221
rect 730 218 782 221
rect 850 218 902 221
rect 906 218 1006 221
rect 1010 218 1030 221
rect 570 208 894 211
rect 1026 208 1134 211
rect 440 203 442 207
rect 446 203 449 207
rect 454 203 456 207
rect 1134 202 1137 208
rect 538 198 638 201
rect 642 198 662 201
rect 666 198 798 201
rect 802 198 846 201
rect 858 198 926 201
rect 962 198 1014 201
rect 1242 198 1302 201
rect 1346 198 1374 201
rect 322 188 350 191
rect 354 188 374 191
rect 450 188 734 191
rect 770 188 1241 191
rect 1238 182 1241 188
rect 402 178 510 181
rect 562 178 686 181
rect 930 178 1118 181
rect 1122 178 1150 181
rect 1154 178 1198 181
rect 1218 178 1230 181
rect 366 171 369 178
rect 366 168 438 171
rect 242 158 310 161
rect 314 158 422 161
rect 510 161 513 168
rect 426 158 513 161
rect 914 158 934 161
rect 954 158 958 161
rect 966 161 969 168
rect 966 158 1118 161
rect 1130 158 1182 161
rect 1198 161 1201 168
rect 1214 161 1217 168
rect 1198 158 1217 161
rect 298 148 374 151
rect 394 148 462 151
rect 474 148 478 151
rect 610 148 638 151
rect 646 148 654 151
rect 658 148 670 151
rect 722 148 734 151
rect 866 148 897 151
rect 922 148 926 151
rect 954 148 1030 151
rect 1034 148 1062 151
rect 1066 148 1254 151
rect 142 142 145 148
rect 894 142 897 148
rect 1358 142 1361 148
rect -26 141 -22 142
rect -26 138 6 141
rect 10 138 14 141
rect 18 138 30 141
rect 410 138 486 141
rect 594 138 694 141
rect 698 138 862 141
rect 930 138 966 141
rect 1018 138 1054 141
rect 1058 138 1134 141
rect 1138 138 1206 141
rect 1210 138 1214 141
rect 406 131 409 138
rect 90 128 161 131
rect 406 128 414 131
rect 550 131 553 138
rect 482 128 553 131
rect 786 128 910 131
rect 938 128 950 131
rect 1018 128 1046 131
rect 1050 128 1078 131
rect 1114 128 1142 131
rect 158 122 161 128
rect 430 121 433 128
rect 378 118 433 121
rect 498 118 614 121
rect 986 118 1030 121
rect 1258 118 1422 121
rect 1426 118 1438 121
rect 986 108 1238 111
rect 1242 108 1342 111
rect 1370 108 1406 111
rect 960 103 962 107
rect 966 103 969 107
rect 974 103 976 107
rect 162 98 182 101
rect 202 98 222 101
rect 330 98 502 101
rect 586 98 854 101
rect 1082 98 1142 101
rect 1242 98 1326 101
rect 322 88 398 91
rect 426 88 486 91
rect 562 88 622 91
rect 818 88 982 91
rect 290 78 350 81
rect 458 78 478 81
rect 522 78 542 81
rect 562 78 590 81
rect 646 81 649 88
rect 646 78 702 81
rect 930 78 958 81
rect 1086 81 1089 88
rect 1334 82 1337 88
rect 1086 78 1118 81
rect 166 71 169 78
rect 166 68 294 71
rect 362 68 430 71
rect 490 68 518 71
rect 698 68 734 71
rect 882 68 990 71
rect 1082 68 1086 71
rect 1114 68 1126 71
rect 298 58 302 61
rect 362 58 366 61
rect 394 58 406 61
rect 474 58 558 61
rect 574 61 577 68
rect 574 58 606 61
rect 642 58 718 61
rect 722 58 726 61
rect 914 58 950 61
rect 1106 58 1254 61
rect 402 48 406 51
rect 498 48 686 51
rect 690 48 702 51
rect 946 48 974 51
rect 986 48 1097 51
rect 1470 51 1474 52
rect 1362 48 1474 51
rect 1094 42 1097 48
rect 538 38 566 41
rect 570 38 646 41
rect 1422 12 1425 18
rect 882 8 1310 11
rect 1314 8 1334 11
rect 1394 8 1406 11
rect 440 3 442 7
rect 446 3 449 7
rect 454 3 456 7
<< m4contact >>
rect 962 1303 966 1307
rect 970 1303 973 1307
rect 973 1303 974 1307
rect 1006 1298 1010 1302
rect 1270 1298 1274 1302
rect 1286 1298 1290 1302
rect 1358 1298 1362 1302
rect 1382 1298 1386 1302
rect 1390 1298 1394 1302
rect 1406 1298 1410 1302
rect 1422 1298 1426 1302
rect 1438 1298 1442 1302
rect 1214 1288 1218 1292
rect 1262 1288 1266 1292
rect 1326 1288 1330 1292
rect 1342 1288 1346 1292
rect 1422 1288 1426 1292
rect 1262 1278 1266 1282
rect 478 1258 482 1262
rect 710 1258 714 1262
rect 1430 1258 1434 1262
rect 286 1248 290 1252
rect 14 1218 18 1222
rect 442 1203 446 1207
rect 450 1203 453 1207
rect 453 1203 454 1207
rect 1406 1198 1410 1202
rect 750 1178 754 1182
rect 1422 1168 1426 1172
rect 1422 1158 1426 1162
rect 862 1148 866 1152
rect 1438 1118 1442 1122
rect 574 1108 578 1112
rect 886 1108 890 1112
rect 998 1108 1002 1112
rect 962 1103 966 1107
rect 970 1103 973 1107
rect 973 1103 974 1107
rect 830 1098 834 1102
rect 742 1078 746 1082
rect 1414 1078 1418 1082
rect 494 1068 498 1072
rect 870 1068 874 1072
rect 878 1068 882 1072
rect 958 1058 962 1062
rect 1102 1058 1106 1062
rect 494 1048 498 1052
rect 878 1048 882 1052
rect 1126 1048 1130 1052
rect 478 1038 482 1042
rect 694 1028 698 1032
rect 742 1028 746 1032
rect 1166 1028 1170 1032
rect 958 1018 962 1022
rect 1430 1008 1434 1012
rect 442 1003 446 1007
rect 450 1003 453 1007
rect 453 1003 454 1007
rect 606 988 610 992
rect 878 988 882 992
rect 1166 988 1170 992
rect 1438 978 1442 982
rect 574 958 578 962
rect 486 948 490 952
rect 766 948 770 952
rect 982 948 986 952
rect 110 938 114 942
rect 750 938 754 942
rect 854 938 858 942
rect 278 918 282 922
rect 462 918 466 922
rect 862 918 866 922
rect 1230 918 1234 922
rect 838 908 842 912
rect 846 908 850 912
rect 962 903 966 907
rect 970 903 973 907
rect 973 903 974 907
rect 14 888 18 892
rect 750 888 754 892
rect 1166 878 1170 882
rect 862 868 866 872
rect 1158 868 1162 872
rect 1238 868 1242 872
rect 110 858 114 862
rect 1334 858 1338 862
rect 854 848 858 852
rect 1102 828 1106 832
rect 486 818 490 822
rect 1126 818 1130 822
rect 442 803 446 807
rect 450 803 453 807
rect 453 803 454 807
rect 846 788 850 792
rect 782 768 786 772
rect 878 768 882 772
rect 942 768 946 772
rect 526 758 530 762
rect 726 758 730 762
rect 782 758 786 762
rect 614 748 618 752
rect 694 748 698 752
rect 718 748 722 752
rect 910 738 914 742
rect 998 738 1002 742
rect 742 718 746 722
rect 862 718 866 722
rect 710 708 714 712
rect 814 708 818 712
rect 962 703 966 707
rect 970 703 973 707
rect 973 703 974 707
rect 526 698 530 702
rect 462 678 466 682
rect 502 678 506 682
rect 894 678 898 682
rect 934 678 938 682
rect 798 668 802 672
rect 942 668 946 672
rect 950 668 954 672
rect 718 658 722 662
rect 726 648 730 652
rect 694 638 698 642
rect 1190 638 1194 642
rect 462 618 466 622
rect 742 608 746 612
rect 442 603 446 607
rect 450 603 453 607
rect 453 603 454 607
rect 870 598 874 602
rect 998 588 1002 592
rect 702 568 706 572
rect 462 558 466 562
rect 774 558 778 562
rect 502 548 506 552
rect 86 528 90 532
rect 782 528 786 532
rect 790 528 794 532
rect 1118 528 1122 532
rect 894 508 898 512
rect 962 503 966 507
rect 970 503 973 507
rect 973 503 974 507
rect 934 498 938 502
rect 1358 498 1362 502
rect 694 488 698 492
rect 798 488 802 492
rect 886 488 890 492
rect 6 478 10 482
rect 638 478 642 482
rect 918 478 922 482
rect 830 468 834 472
rect 902 458 906 462
rect 750 448 754 452
rect 1422 448 1426 452
rect 790 438 794 442
rect 726 428 730 432
rect 442 403 446 407
rect 450 403 453 407
rect 453 403 454 407
rect 1118 398 1122 402
rect 814 388 818 392
rect 782 368 786 372
rect 798 358 802 362
rect 910 358 914 362
rect 918 358 922 362
rect 1198 358 1202 362
rect 1422 358 1426 362
rect 694 348 698 352
rect 774 348 778 352
rect 1214 348 1218 352
rect 1358 348 1362 352
rect 1390 348 1394 352
rect 102 338 106 342
rect 278 338 282 342
rect 718 338 722 342
rect 814 338 818 342
rect 1134 338 1138 342
rect 1414 338 1418 342
rect 542 328 546 332
rect 638 328 642 332
rect 782 328 786 332
rect 494 318 498 322
rect 734 318 738 322
rect 86 308 90 312
rect 502 308 506 312
rect 926 308 930 312
rect 1230 308 1234 312
rect 962 303 966 307
rect 970 303 973 307
rect 973 303 974 307
rect 702 298 706 302
rect 790 298 794 302
rect 830 298 834 302
rect 846 298 850 302
rect 822 278 826 282
rect 70 268 74 272
rect 622 268 626 272
rect 862 268 866 272
rect 1118 268 1122 272
rect 534 258 538 262
rect 822 258 826 262
rect 534 238 538 242
rect 718 238 722 242
rect 750 228 754 232
rect 566 218 570 222
rect 782 218 786 222
rect 566 208 570 212
rect 1134 208 1138 212
rect 442 203 446 207
rect 450 203 453 207
rect 453 203 454 207
rect 846 198 850 202
rect 766 188 770 192
rect 398 178 402 182
rect 950 158 954 162
rect 1118 158 1122 162
rect 470 148 474 152
rect 6 138 10 142
rect 142 138 146 142
rect 694 138 698 142
rect 1206 138 1210 142
rect 1358 138 1362 142
rect 782 128 786 132
rect 950 128 954 132
rect 982 118 986 122
rect 982 108 986 112
rect 1406 108 1410 112
rect 962 103 966 107
rect 970 103 973 107
rect 973 103 974 107
rect 1238 98 1242 102
rect 982 88 986 92
rect 558 78 562 82
rect 1334 78 1338 82
rect 1078 68 1082 72
rect 294 58 298 62
rect 358 58 362 62
rect 726 58 730 62
rect 398 48 402 52
rect 494 48 498 52
rect 702 48 706 52
rect 566 38 570 42
rect 1422 18 1426 22
rect 878 8 882 12
rect 1390 8 1394 12
rect 442 3 446 7
rect 450 3 453 7
rect 453 3 454 7
<< metal4 >>
rect 1270 1308 1345 1311
rect 960 1303 962 1307
rect 966 1303 969 1307
rect 974 1303 976 1307
rect 1270 1302 1273 1308
rect 998 1298 1006 1301
rect 1290 1298 1294 1301
rect 1342 1301 1345 1308
rect 1342 1298 1358 1301
rect 1374 1298 1382 1301
rect 1394 1298 1401 1301
rect 1410 1298 1417 1301
rect 1426 1298 1430 1301
rect 278 1248 286 1251
rect 14 892 17 1218
rect 110 862 113 938
rect 278 922 281 1248
rect 440 1203 442 1207
rect 446 1203 449 1207
rect 454 1203 456 1207
rect 478 1042 481 1258
rect 494 1052 497 1068
rect 440 1003 442 1007
rect 446 1003 449 1007
rect 454 1003 456 1007
rect 574 962 577 1108
rect 698 1028 705 1031
rect 440 803 442 807
rect 446 803 449 807
rect 454 803 456 807
rect 462 682 465 918
rect 486 822 489 948
rect 526 702 529 758
rect 606 751 609 988
rect 606 748 614 751
rect 440 603 442 607
rect 446 603 449 607
rect 454 603 456 607
rect 462 562 465 618
rect 502 552 505 678
rect 694 642 697 748
rect 702 572 705 1028
rect 710 712 713 1258
rect 742 1072 745 1078
rect 742 891 745 1028
rect 750 942 753 1178
rect 834 1098 841 1101
rect 742 888 750 891
rect 718 662 721 748
rect 6 142 9 478
rect 86 312 89 528
rect 440 403 442 407
rect 446 403 449 407
rect 454 403 456 407
rect 278 342 281 348
rect 106 338 110 341
rect 542 332 545 338
rect 638 332 641 478
rect 694 352 697 488
rect 74 268 78 271
rect 440 203 442 207
rect 446 203 449 207
rect 454 203 456 207
rect 146 138 150 141
rect 358 62 361 78
rect 298 58 302 61
rect 398 52 401 178
rect 470 142 473 148
rect 494 52 497 318
rect 502 62 505 308
rect 618 268 622 271
rect 534 242 537 258
rect 566 212 569 218
rect 554 78 558 81
rect 566 42 569 208
rect 694 142 697 348
rect 718 342 721 658
rect 726 652 729 758
rect 742 612 745 718
rect 730 428 737 431
rect 734 322 737 428
rect 702 302 705 308
rect 702 52 705 298
rect 718 61 721 238
rect 750 232 753 448
rect 766 192 769 948
rect 838 912 841 1098
rect 846 792 849 908
rect 854 852 857 938
rect 862 922 865 1148
rect 998 1112 1001 1298
rect 1262 1292 1265 1298
rect 1218 1288 1222 1291
rect 1322 1288 1326 1291
rect 1338 1288 1342 1291
rect 1398 1282 1401 1298
rect 1414 1292 1417 1298
rect 1266 1278 1270 1281
rect 878 1072 881 1078
rect 782 762 785 768
rect 774 352 777 558
rect 782 532 785 758
rect 862 722 865 868
rect 790 442 793 528
rect 798 492 801 668
rect 782 352 785 368
rect 790 361 793 438
rect 814 392 817 708
rect 870 602 873 1068
rect 878 992 881 1048
rect 790 358 798 361
rect 782 222 785 328
rect 790 302 793 358
rect 818 338 825 341
rect 822 282 825 338
rect 830 302 833 468
rect 822 262 825 278
rect 782 132 785 218
rect 846 202 849 298
rect 866 268 870 271
rect 718 58 726 61
rect 878 12 881 768
rect 886 492 889 1108
rect 960 1103 962 1107
rect 966 1103 969 1107
rect 974 1103 976 1107
rect 958 1022 961 1058
rect 960 903 962 907
rect 966 903 969 907
rect 974 903 976 907
rect 898 678 902 681
rect 894 461 897 508
rect 894 458 902 461
rect 910 362 913 738
rect 934 502 937 678
rect 942 672 945 768
rect 960 703 962 707
rect 966 703 969 707
rect 974 703 976 707
rect 950 672 953 678
rect 960 503 962 507
rect 966 503 969 507
rect 974 503 976 507
rect 918 362 921 478
rect 930 308 934 311
rect 934 72 937 308
rect 960 303 962 307
rect 966 303 969 307
rect 974 303 976 307
rect 950 132 953 158
rect 982 122 985 948
rect 1102 832 1105 1058
rect 1126 822 1129 1048
rect 1158 872 1161 1228
rect 1166 992 1169 1028
rect 1166 882 1169 988
rect 998 592 1001 738
rect 1118 402 1121 528
rect 1190 361 1193 638
rect 1190 358 1198 361
rect 1114 268 1118 271
rect 1134 212 1137 338
rect 1118 142 1121 158
rect 1214 141 1217 348
rect 1230 312 1233 918
rect 1210 138 1217 141
rect 960 103 962 107
rect 966 103 969 107
rect 974 103 976 107
rect 982 92 985 108
rect 1238 102 1241 868
rect 1334 82 1337 858
rect 1358 352 1361 498
rect 1354 138 1358 141
rect 1082 68 1086 71
rect 1390 12 1393 348
rect 1406 112 1409 1198
rect 1422 1172 1425 1288
rect 1414 342 1417 1078
rect 1422 452 1425 1158
rect 1430 1012 1433 1258
rect 1438 1232 1441 1298
rect 1438 982 1441 1118
rect 1422 22 1425 358
rect 440 3 442 7
rect 446 3 449 7
rect 454 3 456 7
<< m5contact >>
rect 962 1303 966 1307
rect 969 1303 970 1307
rect 970 1303 973 1307
rect 1262 1298 1266 1302
rect 1294 1298 1298 1302
rect 1382 1298 1386 1302
rect 1430 1298 1434 1302
rect 442 1203 446 1207
rect 449 1203 450 1207
rect 450 1203 453 1207
rect 442 1003 446 1007
rect 449 1003 450 1007
rect 450 1003 453 1007
rect 442 803 446 807
rect 449 803 450 807
rect 450 803 453 807
rect 442 603 446 607
rect 449 603 450 607
rect 450 603 453 607
rect 742 1068 746 1072
rect 442 403 446 407
rect 449 403 450 407
rect 450 403 453 407
rect 278 348 282 352
rect 110 338 114 342
rect 542 338 546 342
rect 78 268 82 272
rect 442 203 446 207
rect 449 203 450 207
rect 450 203 453 207
rect 150 138 154 142
rect 358 78 362 82
rect 302 58 306 62
rect 470 138 474 142
rect 614 268 618 272
rect 550 78 554 82
rect 502 58 506 62
rect 702 308 706 312
rect 1222 1288 1226 1292
rect 1318 1288 1322 1292
rect 1334 1288 1338 1292
rect 1414 1288 1418 1292
rect 1270 1278 1274 1282
rect 1398 1278 1402 1282
rect 1158 1228 1162 1232
rect 878 1078 882 1082
rect 782 348 786 352
rect 870 268 874 272
rect 962 1103 966 1107
rect 969 1103 970 1107
rect 970 1103 973 1107
rect 962 903 966 907
rect 969 903 970 907
rect 970 903 973 907
rect 902 678 906 682
rect 962 703 966 707
rect 969 703 970 707
rect 970 703 973 707
rect 950 678 954 682
rect 962 503 966 507
rect 969 503 970 507
rect 970 503 973 507
rect 934 308 938 312
rect 962 303 966 307
rect 969 303 970 307
rect 970 303 973 307
rect 1110 268 1114 272
rect 1118 138 1122 142
rect 962 103 966 107
rect 969 103 970 107
rect 970 103 973 107
rect 1350 138 1354 142
rect 934 68 938 72
rect 1086 68 1090 72
rect 1438 1228 1442 1232
rect 442 3 446 7
rect 449 3 450 7
rect 450 3 453 7
<< metal5 >>
rect 966 1303 969 1307
rect 965 1302 970 1303
rect 975 1302 976 1307
rect 1266 1298 1277 1301
rect 1298 1298 1377 1301
rect 1386 1298 1430 1301
rect 1226 1288 1318 1291
rect 1330 1288 1334 1291
rect 1374 1291 1377 1298
rect 1374 1288 1414 1291
rect 1274 1278 1398 1281
rect 1162 1228 1438 1231
rect 446 1203 449 1207
rect 445 1202 450 1203
rect 455 1202 456 1207
rect 966 1103 969 1107
rect 965 1102 970 1103
rect 975 1102 976 1107
rect 878 1071 881 1078
rect 746 1068 881 1071
rect 446 1003 449 1007
rect 445 1002 450 1003
rect 455 1002 456 1007
rect 966 903 969 907
rect 965 902 970 903
rect 975 902 976 907
rect 446 803 449 807
rect 445 802 450 803
rect 455 802 456 807
rect 966 703 969 707
rect 965 702 970 703
rect 975 702 976 707
rect 906 678 950 681
rect 446 603 449 607
rect 445 602 450 603
rect 455 602 456 607
rect 966 503 969 507
rect 965 502 970 503
rect 975 502 976 507
rect 446 403 449 407
rect 445 402 450 403
rect 455 402 456 407
rect 282 348 782 351
rect 114 338 542 341
rect 706 308 934 311
rect 966 303 969 307
rect 965 302 970 303
rect 975 302 976 307
rect 82 268 614 271
rect 874 268 1110 271
rect 446 203 449 207
rect 445 202 450 203
rect 455 202 456 207
rect 154 138 470 141
rect 1122 138 1350 141
rect 966 103 969 107
rect 965 102 970 103
rect 975 102 976 107
rect 362 78 550 81
rect 938 68 1086 71
rect 306 58 502 61
rect 446 3 449 7
rect 445 2 450 3
rect 455 2 456 7
<< m6contact >>
rect 960 1303 962 1307
rect 962 1303 965 1307
rect 970 1303 973 1307
rect 973 1303 975 1307
rect 960 1302 965 1303
rect 970 1302 975 1303
rect 1277 1297 1282 1302
rect 1325 1287 1330 1292
rect 440 1203 442 1207
rect 442 1203 445 1207
rect 450 1203 453 1207
rect 453 1203 455 1207
rect 440 1202 445 1203
rect 450 1202 455 1203
rect 960 1103 962 1107
rect 962 1103 965 1107
rect 970 1103 973 1107
rect 973 1103 975 1107
rect 960 1102 965 1103
rect 970 1102 975 1103
rect 440 1003 442 1007
rect 442 1003 445 1007
rect 450 1003 453 1007
rect 453 1003 455 1007
rect 440 1002 445 1003
rect 450 1002 455 1003
rect 960 903 962 907
rect 962 903 965 907
rect 970 903 973 907
rect 973 903 975 907
rect 960 902 965 903
rect 970 902 975 903
rect 440 803 442 807
rect 442 803 445 807
rect 450 803 453 807
rect 453 803 455 807
rect 440 802 445 803
rect 450 802 455 803
rect 960 703 962 707
rect 962 703 965 707
rect 970 703 973 707
rect 973 703 975 707
rect 960 702 965 703
rect 970 702 975 703
rect 440 603 442 607
rect 442 603 445 607
rect 450 603 453 607
rect 453 603 455 607
rect 440 602 445 603
rect 450 602 455 603
rect 960 503 962 507
rect 962 503 965 507
rect 970 503 973 507
rect 973 503 975 507
rect 960 502 965 503
rect 970 502 975 503
rect 440 403 442 407
rect 442 403 445 407
rect 450 403 453 407
rect 453 403 455 407
rect 440 402 445 403
rect 450 402 455 403
rect 960 303 962 307
rect 962 303 965 307
rect 970 303 973 307
rect 973 303 975 307
rect 960 302 965 303
rect 970 302 975 303
rect 440 203 442 207
rect 442 203 445 207
rect 450 203 453 207
rect 453 203 455 207
rect 440 202 445 203
rect 450 202 455 203
rect 960 103 962 107
rect 962 103 965 107
rect 970 103 973 107
rect 973 103 975 107
rect 960 102 965 103
rect 970 102 975 103
rect 440 3 442 7
rect 442 3 445 7
rect 450 3 453 7
rect 453 3 455 7
rect 440 2 445 3
rect 450 2 455 3
<< metal6 >>
rect 440 1207 456 1330
rect 445 1202 450 1207
rect 455 1202 456 1207
rect 440 1007 456 1202
rect 445 1002 450 1007
rect 455 1002 456 1007
rect 440 807 456 1002
rect 445 802 450 807
rect 455 802 456 807
rect 440 607 456 802
rect 445 602 450 607
rect 455 602 456 607
rect 440 407 456 602
rect 445 402 450 407
rect 455 402 456 407
rect 440 207 456 402
rect 445 202 450 207
rect 455 202 456 207
rect 440 7 456 202
rect 445 2 450 7
rect 455 2 456 7
rect 440 -30 456 2
rect 960 1307 976 1330
rect 965 1302 970 1307
rect 975 1302 976 1307
rect 960 1107 976 1302
rect 1277 1307 1330 1312
rect 1277 1302 1282 1307
rect 1325 1292 1330 1307
rect 965 1102 970 1107
rect 975 1102 976 1107
rect 960 907 976 1102
rect 965 902 970 907
rect 975 902 976 907
rect 960 707 976 902
rect 965 702 970 707
rect 975 702 976 707
rect 960 507 976 702
rect 965 502 970 507
rect 975 502 976 507
rect 960 307 976 502
rect 965 302 970 307
rect 975 302 976 307
rect 960 107 976 302
rect 965 102 970 107
rect 975 102 976 107
rect 960 -30 976 102
use PADFC  PADFC_0
timestamp 1560662619
transform 1 0 -3098 0 1 1536
box 0 0 3000 3000
use PADVDD  PADVDD_0
timestamp 1560662619
transform 1 0 -98 0 1 1536
box 0 0 900 3000
use PADVDD  PADVDD_1
timestamp 1560662619
transform 1 0 802 0 1 1536
box 0 0 900 3000
use PADFC  PADFC_1
timestamp 1560662619
transform 0 1 1666 -1 0 4536
box 0 0 3000 3000
use PADINC  PADINC_2
timestamp 1560662619
transform 0 -1 -98 1 0 648
box 0 0 900 3000
use INVX8  INVX8_4
timestamp 1560662619
transform 1 0 4 0 -1 1305
box 0 0 40 100
use INVX8  INVX8_1
timestamp 1560662619
transform 1 0 44 0 -1 1305
box 0 0 40 100
use DFFSR  DFFSR_32
timestamp 1560662619
transform -1 0 260 0 -1 1305
box 0 0 176 100
use BUFX2  BUFX2_24
timestamp 1560662619
transform -1 0 284 0 -1 1305
box 0 0 24 100
use DFFSR  DFFSR_28
timestamp 1560662619
transform 1 0 284 0 -1 1305
box 0 0 176 100
use FILL  FILL_12_0_0
timestamp 1560662619
transform 1 0 460 0 -1 1305
box 0 0 8 100
use FILL  FILL_12_0_1
timestamp 1560662619
transform 1 0 468 0 -1 1305
box 0 0 8 100
use BUFX2  BUFX2_23
timestamp 1560662619
transform 1 0 476 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_38
timestamp 1560662619
transform -1 0 524 0 -1 1305
box 0 0 24 100
use DFFSR  DFFSR_31
timestamp 1560662619
transform -1 0 700 0 -1 1305
box 0 0 176 100
use BUFX4  BUFX4_6
timestamp 1560662619
transform -1 0 732 0 -1 1305
box 0 0 32 100
use INVX1  INVX1_12
timestamp 1560662619
transform 1 0 732 0 -1 1305
box 0 0 16 100
use DFFSR  DFFSR_1
timestamp 1560662619
transform -1 0 924 0 -1 1305
box 0 0 176 100
use BUFX2  BUFX2_22
timestamp 1560662619
transform -1 0 948 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_35
timestamp 1560662619
transform 1 0 948 0 -1 1305
box 0 0 24 100
use FILL  FILL_12_1_0
timestamp 1560662619
transform -1 0 980 0 -1 1305
box 0 0 8 100
use FILL  FILL_12_1_1
timestamp 1560662619
transform -1 0 988 0 -1 1305
box 0 0 8 100
use DFFSR  DFFSR_5
timestamp 1560662619
transform -1 0 1164 0 -1 1305
box 0 0 176 100
use BUFX2  BUFX2_29
timestamp 1560662619
transform 1 0 1164 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_30
timestamp 1560662619
transform 1 0 1188 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_32
timestamp 1560662619
transform 1 0 1212 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_31
timestamp 1560662619
transform 1 0 1236 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_33
timestamp 1560662619
transform 1 0 1260 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_27
timestamp 1560662619
transform 1 0 1284 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_28
timestamp 1560662619
transform 1 0 1308 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_17
timestamp 1560662619
transform 1 0 1332 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_34
timestamp 1560662619
transform 1 0 1356 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_15
timestamp 1560662619
transform 1 0 1380 0 -1 1305
box 0 0 24 100
use BUFX2  BUFX2_18
timestamp 1560662619
transform 1 0 1404 0 -1 1305
box 0 0 24 100
use FILL  FILL_13_1
timestamp 1560662619
transform -1 0 1436 0 -1 1305
box 0 0 8 100
use FILL  FILL_13_2
timestamp 1560662619
transform -1 0 1444 0 -1 1305
box 0 0 8 100
use BUFX2  BUFX2_37
timestamp 1560662619
transform -1 0 28 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_1
timestamp 1560662619
transform -1 0 52 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_25
timestamp 1560662619
transform 1 0 52 0 1 1105
box 0 0 24 100
use DFFSR  DFFSR_24
timestamp 1560662619
transform -1 0 252 0 1 1105
box 0 0 176 100
use NAND2X1  NAND2X1_45
timestamp 1560662619
transform 1 0 252 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_49
timestamp 1560662619
transform -1 0 308 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_48
timestamp 1560662619
transform -1 0 340 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_41
timestamp 1560662619
transform 1 0 340 0 1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_41
timestamp 1560662619
transform -1 0 396 0 1 1105
box 0 0 24 100
use FILL  FILL_11_0_0
timestamp 1560662619
transform 1 0 396 0 1 1105
box 0 0 8 100
use FILL  FILL_11_0_1
timestamp 1560662619
transform 1 0 404 0 1 1105
box 0 0 8 100
use DFFSR  DFFSR_30
timestamp 1560662619
transform 1 0 412 0 1 1105
box 0 0 176 100
use NAND2X1  NAND2X1_44
timestamp 1560662619
transform 1 0 588 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_47
timestamp 1560662619
transform -1 0 644 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_46
timestamp 1560662619
transform -1 0 676 0 1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_43
timestamp 1560662619
transform 1 0 676 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_45
timestamp 1560662619
transform -1 0 732 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_42
timestamp 1560662619
transform 1 0 732 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_44
timestamp 1560662619
transform -1 0 796 0 1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_43
timestamp 1560662619
transform 1 0 796 0 1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_42
timestamp 1560662619
transform -1 0 852 0 1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_5
timestamp 1560662619
transform 1 0 852 0 1 1105
box 0 0 48 100
use FILL  FILL_11_1_0
timestamp 1560662619
transform -1 0 908 0 1 1105
box 0 0 8 100
use FILL  FILL_11_1_1
timestamp 1560662619
transform -1 0 916 0 1 1105
box 0 0 8 100
use DFFSR  DFFSR_29
timestamp 1560662619
transform -1 0 1092 0 1 1105
box 0 0 176 100
use INVX1  INVX1_22
timestamp 1560662619
transform 1 0 1092 0 1 1105
box 0 0 16 100
use AOI21X1  AOI21X1_4
timestamp 1560662619
transform 1 0 1108 0 1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_15
timestamp 1560662619
transform -1 0 1164 0 1 1105
box 0 0 24 100
use DFFSR  DFFSR_2
timestamp 1560662619
transform -1 0 1340 0 1 1105
box 0 0 176 100
use BUFX2  BUFX2_26
timestamp 1560662619
transform 1 0 1340 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_11
timestamp 1560662619
transform 1 0 1364 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_13
timestamp 1560662619
transform 1 0 1388 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_9
timestamp 1560662619
transform 1 0 1412 0 1 1105
box 0 0 24 100
use FILL  FILL_12_1
timestamp 1560662619
transform 1 0 1436 0 1 1105
box 0 0 8 100
use INVX1  INVX1_8
timestamp 1560662619
transform -1 0 20 0 -1 1105
box 0 0 16 100
use DFFSR  DFFSR_27
timestamp 1560662619
transform 1 0 20 0 -1 1105
box 0 0 176 100
use NAND2X1  NAND2X1_40
timestamp 1560662619
transform 1 0 196 0 -1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_39
timestamp 1560662619
transform -1 0 252 0 -1 1105
box 0 0 32 100
use INVX4  INVX4_4
timestamp 1560662619
transform -1 0 276 0 -1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_38
timestamp 1560662619
transform -1 0 308 0 -1 1105
box 0 0 32 100
use OAI21X1  OAI21X1_40
timestamp 1560662619
transform 1 0 308 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_39
timestamp 1560662619
transform 1 0 340 0 -1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_37
timestamp 1560662619
transform -1 0 396 0 -1 1105
box 0 0 32 100
use FILL  FILL_10_0_0
timestamp 1560662619
transform -1 0 404 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_0_1
timestamp 1560662619
transform -1 0 412 0 -1 1105
box 0 0 8 100
use DFFSR  DFFSR_26
timestamp 1560662619
transform -1 0 588 0 -1 1105
box 0 0 176 100
use OAI21X1  OAI21X1_36
timestamp 1560662619
transform -1 0 620 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_44
timestamp 1560662619
transform -1 0 644 0 -1 1105
box 0 0 24 100
use INVX1  INVX1_38
timestamp 1560662619
transform 1 0 644 0 -1 1105
box 0 0 16 100
use OAI21X1  OAI21X1_35
timestamp 1560662619
transform 1 0 660 0 -1 1105
box 0 0 32 100
use NAND3X1  NAND3X1_20
timestamp 1560662619
transform -1 0 724 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_43
timestamp 1560662619
transform -1 0 748 0 -1 1105
box 0 0 24 100
use NOR2X1  NOR2X1_42
timestamp 1560662619
transform -1 0 772 0 -1 1105
box 0 0 24 100
use DFFSR  DFFSR_25
timestamp 1560662619
transform -1 0 948 0 -1 1105
box 0 0 176 100
use NAND2X1  NAND2X1_12
timestamp 1560662619
transform -1 0 972 0 -1 1105
box 0 0 24 100
use FILL  FILL_10_1_0
timestamp 1560662619
transform 1 0 972 0 -1 1105
box 0 0 8 100
use FILL  FILL_10_1_1
timestamp 1560662619
transform 1 0 980 0 -1 1105
box 0 0 8 100
use BUFX2  BUFX2_21
timestamp 1560662619
transform 1 0 988 0 -1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_2
timestamp 1560662619
transform 1 0 1012 0 -1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_13
timestamp 1560662619
transform 1 0 1044 0 -1 1105
box 0 0 24 100
use AOI22X1  AOI22X1_1
timestamp 1560662619
transform 1 0 1068 0 -1 1105
box 0 0 40 100
use NAND2X1  NAND2X1_13
timestamp 1560662619
transform 1 0 1108 0 -1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_4
timestamp 1560662619
transform 1 0 1132 0 -1 1105
box 0 0 32 100
use DFFSR  DFFSR_11
timestamp 1560662619
transform 1 0 1164 0 -1 1105
box 0 0 176 100
use BUFX2  BUFX2_36
timestamp 1560662619
transform 1 0 1340 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_7
timestamp 1560662619
transform 1 0 1364 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_2
timestamp 1560662619
transform 1 0 1388 0 -1 1105
box 0 0 24 100
use BUFX2  BUFX2_8
timestamp 1560662619
transform 1 0 1412 0 -1 1105
box 0 0 24 100
use FILL  FILL_11_1
timestamp 1560662619
transform -1 0 1444 0 -1 1105
box 0 0 8 100
use DFFSR  DFFSR_8
timestamp 1560662619
transform -1 0 180 0 1 905
box 0 0 176 100
use DFFSR  DFFSR_7
timestamp 1560662619
transform 1 0 180 0 1 905
box 0 0 176 100
use NOR2X1  NOR2X1_41
timestamp 1560662619
transform 1 0 356 0 1 905
box 0 0 24 100
use NOR2X1  NOR2X1_40
timestamp 1560662619
transform 1 0 380 0 1 905
box 0 0 24 100
use NOR2X1  NOR2X1_39
timestamp 1560662619
transform -1 0 428 0 1 905
box 0 0 24 100
use INVX4  INVX4_3
timestamp 1560662619
transform 1 0 428 0 1 905
box 0 0 24 100
use FILL  FILL_9_0_0
timestamp 1560662619
transform 1 0 452 0 1 905
box 0 0 8 100
use FILL  FILL_9_0_1
timestamp 1560662619
transform 1 0 460 0 1 905
box 0 0 8 100
use INVX1  INVX1_16
timestamp 1560662619
transform 1 0 468 0 1 905
box 0 0 16 100
use AOI21X1  AOI21X1_3
timestamp 1560662619
transform 1 0 484 0 1 905
box 0 0 32 100
use NOR2X1  NOR2X1_14
timestamp 1560662619
transform -1 0 540 0 1 905
box 0 0 24 100
use DFFSR  DFFSR_4
timestamp 1560662619
transform 1 0 540 0 1 905
box 0 0 176 100
use NOR2X1  NOR2X1_45
timestamp 1560662619
transform -1 0 740 0 1 905
box 0 0 24 100
use OAI22X1  OAI22X1_2
timestamp 1560662619
transform -1 0 780 0 1 905
box 0 0 40 100
use OAI22X1  OAI22X1_1
timestamp 1560662619
transform 1 0 780 0 1 905
box 0 0 40 100
use NAND3X1  NAND3X1_7
timestamp 1560662619
transform 1 0 820 0 1 905
box 0 0 32 100
use NAND3X1  NAND3X1_5
timestamp 1560662619
transform 1 0 852 0 1 905
box 0 0 32 100
use NAND2X1  NAND2X1_10
timestamp 1560662619
transform -1 0 908 0 1 905
box 0 0 24 100
use INVX1  INVX1_21
timestamp 1560662619
transform 1 0 908 0 1 905
box 0 0 16 100
use MUX2X1  MUX2X1_4
timestamp 1560662619
transform -1 0 972 0 1 905
box 0 0 48 100
use FILL  FILL_9_1_0
timestamp 1560662619
transform -1 0 980 0 1 905
box 0 0 8 100
use FILL  FILL_9_1_1
timestamp 1560662619
transform -1 0 988 0 1 905
box 0 0 8 100
use INVX1  INVX1_13
timestamp 1560662619
transform -1 0 1004 0 1 905
box 0 0 16 100
use AOI21X1  AOI21X1_1
timestamp 1560662619
transform -1 0 1036 0 1 905
box 0 0 32 100
use NAND3X1  NAND3X1_2
timestamp 1560662619
transform -1 0 1068 0 1 905
box 0 0 32 100
use DFFSR  DFFSR_3
timestamp 1560662619
transform 1 0 1068 0 1 905
box 0 0 176 100
use DFFSR  DFFSR_10
timestamp 1560662619
transform 1 0 1244 0 1 905
box 0 0 176 100
use BUFX2  BUFX2_20
timestamp 1560662619
transform 1 0 1420 0 1 905
box 0 0 24 100
use BUFX4  BUFX4_10
timestamp 1560662619
transform 1 0 4 0 -1 905
box 0 0 32 100
use DFFSR  DFFSR_21
timestamp 1560662619
transform 1 0 36 0 -1 905
box 0 0 176 100
use INVX1  INVX1_31
timestamp 1560662619
transform 1 0 212 0 -1 905
box 0 0 16 100
use INVX1  INVX1_18
timestamp 1560662619
transform 1 0 228 0 -1 905
box 0 0 16 100
use MUX2X1  MUX2X1_2
timestamp 1560662619
transform -1 0 292 0 -1 905
box 0 0 48 100
use INVX1  INVX1_7
timestamp 1560662619
transform -1 0 308 0 -1 905
box 0 0 16 100
use NOR2X1  NOR2X1_9
timestamp 1560662619
transform 1 0 308 0 -1 905
box 0 0 24 100
use OAI21X1  OAI21X1_3
timestamp 1560662619
transform 1 0 332 0 -1 905
box 0 0 32 100
use INVX1  INVX1_5
timestamp 1560662619
transform -1 0 380 0 -1 905
box 0 0 16 100
use FILL  FILL_8_0_0
timestamp 1560662619
transform -1 0 388 0 -1 905
box 0 0 8 100
use FILL  FILL_8_0_1
timestamp 1560662619
transform -1 0 396 0 -1 905
box 0 0 8 100
use DFFSR  DFFSR_17
timestamp 1560662619
transform -1 0 572 0 -1 905
box 0 0 176 100
use DFFSR  DFFSR_16
timestamp 1560662619
transform 1 0 572 0 -1 905
box 0 0 176 100
use NAND2X1  NAND2X1_11
timestamp 1560662619
transform 1 0 748 0 -1 905
box 0 0 24 100
use INVX4  INVX4_1
timestamp 1560662619
transform -1 0 796 0 -1 905
box 0 0 24 100
use NOR2X1  NOR2X1_4
timestamp 1560662619
transform 1 0 796 0 -1 905
box 0 0 24 100
use NOR3X1  NOR3X1_7
timestamp 1560662619
transform -1 0 884 0 -1 905
box 0 0 64 100
use INVX1  INVX1_2
timestamp 1560662619
transform 1 0 884 0 -1 905
box 0 0 16 100
use NAND2X1  NAND2X1_5
timestamp 1560662619
transform 1 0 900 0 -1 905
box 0 0 24 100
use NOR2X1  NOR2X1_12
timestamp 1560662619
transform -1 0 948 0 -1 905
box 0 0 24 100
use FILL  FILL_8_1_0
timestamp 1560662619
transform -1 0 956 0 -1 905
box 0 0 8 100
use FILL  FILL_8_1_1
timestamp 1560662619
transform -1 0 964 0 -1 905
box 0 0 8 100
use NOR3X1  NOR3X1_2
timestamp 1560662619
transform -1 0 1028 0 -1 905
box 0 0 64 100
use NAND2X1  NAND2X1_4
timestamp 1560662619
transform 1 0 1028 0 -1 905
box 0 0 24 100
use NAND2X1  NAND2X1_15
timestamp 1560662619
transform 1 0 1052 0 -1 905
box 0 0 24 100
use NOR3X1  NOR3X1_6
timestamp 1560662619
transform -1 0 1140 0 -1 905
box 0 0 64 100
use NAND2X1  NAND2X1_7
timestamp 1560662619
transform -1 0 1164 0 -1 905
box 0 0 24 100
use INVX1  INVX1_14
timestamp 1560662619
transform 1 0 1164 0 -1 905
box 0 0 16 100
use OAI21X1  OAI21X1_5
timestamp 1560662619
transform -1 0 1212 0 -1 905
box 0 0 32 100
use OAI21X1  OAI21X1_6
timestamp 1560662619
transform -1 0 1244 0 -1 905
box 0 0 32 100
use DFFSR  DFFSR_9
timestamp 1560662619
transform 1 0 1244 0 -1 905
box 0 0 176 100
use BUFX2  BUFX2_12
timestamp 1560662619
transform 1 0 1420 0 -1 905
box 0 0 24 100
use CLKBUF1  CLKBUF1_1
timestamp 1560662619
transform 1 0 4 0 1 705
box 0 0 72 100
use MUX2X1  MUX2X1_3
timestamp 1560662619
transform -1 0 124 0 1 705
box 0 0 48 100
use INVX1  INVX1_19
timestamp 1560662619
transform -1 0 140 0 1 705
box 0 0 16 100
use MUX2X1  MUX2X1_11
timestamp 1560662619
transform -1 0 188 0 1 705
box 0 0 48 100
use INVX1  INVX1_17
timestamp 1560662619
transform 1 0 188 0 1 705
box 0 0 16 100
use MUX2X1  MUX2X1_1
timestamp 1560662619
transform -1 0 252 0 1 705
box 0 0 48 100
use DFFSR  DFFSR_6
timestamp 1560662619
transform 1 0 252 0 1 705
box 0 0 176 100
use OAI21X1  OAI21X1_1
timestamp 1560662619
transform 1 0 428 0 1 705
box 0 0 32 100
use FILL  FILL_7_0_0
timestamp 1560662619
transform -1 0 468 0 1 705
box 0 0 8 100
use FILL  FILL_7_0_1
timestamp 1560662619
transform -1 0 476 0 1 705
box 0 0 8 100
use INVX1  INVX1_20
timestamp 1560662619
transform -1 0 492 0 1 705
box 0 0 16 100
use BUFX4  BUFX4_8
timestamp 1560662619
transform -1 0 524 0 1 705
box 0 0 32 100
use INVX1  INVX1_27
timestamp 1560662619
transform 1 0 524 0 1 705
box 0 0 16 100
use MUX2X1  MUX2X1_7
timestamp 1560662619
transform -1 0 588 0 1 705
box 0 0 48 100
use CLKBUF1  CLKBUF1_4
timestamp 1560662619
transform 1 0 588 0 1 705
box 0 0 72 100
use MUX2X1  MUX2X1_6
timestamp 1560662619
transform -1 0 708 0 1 705
box 0 0 48 100
use INVX1  INVX1_26
timestamp 1560662619
transform -1 0 724 0 1 705
box 0 0 16 100
use OAI21X1  OAI21X1_2
timestamp 1560662619
transform -1 0 756 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_3
timestamp 1560662619
transform -1 0 788 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_5
timestamp 1560662619
transform -1 0 812 0 1 705
box 0 0 24 100
use NAND3X1  NAND3X1_6
timestamp 1560662619
transform -1 0 844 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_4
timestamp 1560662619
transform -1 0 876 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_1
timestamp 1560662619
transform 1 0 876 0 1 705
box 0 0 32 100
use NAND2X1  NAND2X1_2
timestamp 1560662619
transform 1 0 908 0 1 705
box 0 0 24 100
use INVX1  INVX1_1
timestamp 1560662619
transform -1 0 948 0 1 705
box 0 0 16 100
use NAND3X1  NAND3X1_8
timestamp 1560662619
transform -1 0 980 0 1 705
box 0 0 32 100
use FILL  FILL_7_1_0
timestamp 1560662619
transform -1 0 988 0 1 705
box 0 0 8 100
use FILL  FILL_7_1_1
timestamp 1560662619
transform -1 0 996 0 1 705
box 0 0 8 100
use NOR2X1  NOR2X1_11
timestamp 1560662619
transform -1 0 1020 0 1 705
box 0 0 24 100
use NOR3X1  NOR3X1_1
timestamp 1560662619
transform 1 0 1020 0 1 705
box 0 0 64 100
use NAND2X1  NAND2X1_14
timestamp 1560662619
transform 1 0 1084 0 1 705
box 0 0 24 100
use INVX2  INVX2_1
timestamp 1560662619
transform -1 0 1124 0 1 705
box 0 0 16 100
use NAND3X1  NAND3X1_9
timestamp 1560662619
transform -1 0 1156 0 1 705
box 0 0 32 100
use NAND3X1  NAND3X1_10
timestamp 1560662619
transform 1 0 1156 0 1 705
box 0 0 32 100
use NOR3X1  NOR3X1_5
timestamp 1560662619
transform 1 0 1188 0 1 705
box 0 0 64 100
use DFFSR  DFFSR_45
timestamp 1560662619
transform -1 0 1428 0 1 705
box 0 0 176 100
use FILL  FILL_8_1
timestamp 1560662619
transform 1 0 1428 0 1 705
box 0 0 8 100
use FILL  FILL_8_2
timestamp 1560662619
transform 1 0 1436 0 1 705
box 0 0 8 100
use DFFSR  DFFSR_22
timestamp 1560662619
transform 1 0 4 0 -1 705
box 0 0 176 100
use INVX1  INVX1_30
timestamp 1560662619
transform -1 0 196 0 -1 705
box 0 0 16 100
use INVX1  INVX1_32
timestamp 1560662619
transform 1 0 196 0 -1 705
box 0 0 16 100
use MUX2X1  MUX2X1_12
timestamp 1560662619
transform -1 0 260 0 -1 705
box 0 0 48 100
use DFFSR  DFFSR_18
timestamp 1560662619
transform 1 0 260 0 -1 705
box 0 0 176 100
use INVX1  INVX1_29
timestamp 1560662619
transform -1 0 452 0 -1 705
box 0 0 16 100
use FILL  FILL_6_0_0
timestamp 1560662619
transform -1 0 460 0 -1 705
box 0 0 8 100
use FILL  FILL_6_0_1
timestamp 1560662619
transform -1 0 468 0 -1 705
box 0 0 8 100
use MUX2X1  MUX2X1_9
timestamp 1560662619
transform -1 0 516 0 -1 705
box 0 0 48 100
use INVX1  INVX1_28
timestamp 1560662619
transform 1 0 516 0 -1 705
box 0 0 16 100
use MUX2X1  MUX2X1_8
timestamp 1560662619
transform -1 0 580 0 -1 705
box 0 0 48 100
use INVX4  INVX4_5
timestamp 1560662619
transform -1 0 604 0 -1 705
box 0 0 24 100
use OAI21X1  OAI21X1_27
timestamp 1560662619
transform 1 0 604 0 -1 705
box 0 0 32 100
use DFFSR  DFFSR_36
timestamp 1560662619
transform -1 0 812 0 -1 705
box 0 0 176 100
use NAND2X1  NAND2X1_9
timestamp 1560662619
transform -1 0 836 0 -1 705
box 0 0 24 100
use INVX1  INVX1_6
timestamp 1560662619
transform 1 0 836 0 -1 705
box 0 0 16 100
use NOR2X1  NOR2X1_6
timestamp 1560662619
transform 1 0 852 0 -1 705
box 0 0 24 100
use NOR2X1  NOR2X1_10
timestamp 1560662619
transform -1 0 900 0 -1 705
box 0 0 24 100
use NOR2X1  NOR2X1_3
timestamp 1560662619
transform 1 0 900 0 -1 705
box 0 0 24 100
use INVX2  INVX2_9
timestamp 1560662619
transform 1 0 924 0 -1 705
box 0 0 16 100
use NOR2X1  NOR2X1_7
timestamp 1560662619
transform 1 0 940 0 -1 705
box 0 0 24 100
use FILL  FILL_6_1_0
timestamp 1560662619
transform -1 0 972 0 -1 705
box 0 0 8 100
use FILL  FILL_6_1_1
timestamp 1560662619
transform -1 0 980 0 -1 705
box 0 0 8 100
use INVX1  INVX1_3
timestamp 1560662619
transform -1 0 996 0 -1 705
box 0 0 16 100
use NAND2X1  NAND2X1_6
timestamp 1560662619
transform -1 0 1020 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_3
timestamp 1560662619
transform -1 0 1044 0 -1 705
box 0 0 24 100
use INVX1  INVX1_4
timestamp 1560662619
transform 1 0 1044 0 -1 705
box 0 0 16 100
use NOR2X1  NOR2X1_8
timestamp 1560662619
transform -1 0 1084 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_8
timestamp 1560662619
transform 1 0 1084 0 -1 705
box 0 0 24 100
use NOR3X1  NOR3X1_4
timestamp 1560662619
transform 1 0 1108 0 -1 705
box 0 0 64 100
use NOR3X1  NOR3X1_3
timestamp 1560662619
transform 1 0 1172 0 -1 705
box 0 0 64 100
use DFFSR  DFFSR_44
timestamp 1560662619
transform -1 0 1412 0 -1 705
box 0 0 176 100
use BUFX2  BUFX2_6
timestamp 1560662619
transform 1 0 1412 0 -1 705
box 0 0 24 100
use FILL  FILL_7_1
timestamp 1560662619
transform -1 0 1444 0 -1 705
box 0 0 8 100
use DFFSR  DFFSR_20
timestamp 1560662619
transform 1 0 4 0 1 505
box 0 0 176 100
use MUX2X1  MUX2X1_10
timestamp 1560662619
transform -1 0 228 0 1 505
box 0 0 48 100
use DFFSR  DFFSR_19
timestamp 1560662619
transform 1 0 228 0 1 505
box 0 0 176 100
use XNOR2X1  XNOR2X1_2
timestamp 1560662619
transform -1 0 460 0 1 505
box 0 0 56 100
use FILL  FILL_5_0_0
timestamp 1560662619
transform 1 0 460 0 1 505
box 0 0 8 100
use FILL  FILL_5_0_1
timestamp 1560662619
transform 1 0 468 0 1 505
box 0 0 8 100
use DFFSR  DFFSR_47
timestamp 1560662619
transform 1 0 476 0 1 505
box 0 0 176 100
use INVX1  INVX1_23
timestamp 1560662619
transform 1 0 652 0 1 505
box 0 0 16 100
use OAI21X1  OAI21X1_12
timestamp 1560662619
transform 1 0 668 0 1 505
box 0 0 32 100
use OAI21X1  OAI21X1_28
timestamp 1560662619
transform -1 0 732 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_28
timestamp 1560662619
transform -1 0 756 0 1 505
box 0 0 24 100
use NAND2X1  NAND2X1_32
timestamp 1560662619
transform 1 0 756 0 1 505
box 0 0 24 100
use OAI21X1  OAI21X1_10
timestamp 1560662619
transform 1 0 780 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_18
timestamp 1560662619
transform 1 0 812 0 1 505
box 0 0 24 100
use DFFSR  DFFSR_23
timestamp 1560662619
transform 1 0 836 0 1 505
box 0 0 176 100
use FILL  FILL_5_1_0
timestamp 1560662619
transform 1 0 1012 0 1 505
box 0 0 8 100
use FILL  FILL_5_1_1
timestamp 1560662619
transform 1 0 1020 0 1 505
box 0 0 8 100
use NOR2X1  NOR2X1_46
timestamp 1560662619
transform 1 0 1028 0 1 505
box 0 0 24 100
use OAI21X1  OAI21X1_50
timestamp 1560662619
transform -1 0 1084 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_2
timestamp 1560662619
transform -1 0 1116 0 1 505
box 0 0 32 100
use NOR2X1  NOR2X1_26
timestamp 1560662619
transform -1 0 1140 0 1 505
box 0 0 24 100
use NAND3X1  NAND3X1_11
timestamp 1560662619
transform 1 0 1140 0 1 505
box 0 0 32 100
use INVX1  INVX1_9
timestamp 1560662619
transform -1 0 1188 0 1 505
box 0 0 16 100
use DFFSR  DFFSR_46
timestamp 1560662619
transform -1 0 1364 0 1 505
box 0 0 176 100
use CLKBUF1  CLKBUF1_3
timestamp 1560662619
transform -1 0 1436 0 1 505
box 0 0 72 100
use FILL  FILL_6_1
timestamp 1560662619
transform 1 0 1436 0 1 505
box 0 0 8 100
use BUFX4  BUFX4_5
timestamp 1560662619
transform 1 0 4 0 -1 505
box 0 0 32 100
use DFFSR  DFFSR_37
timestamp 1560662619
transform 1 0 36 0 -1 505
box 0 0 176 100
use DFFSR  DFFSR_39
timestamp 1560662619
transform 1 0 212 0 -1 505
box 0 0 176 100
use OAI21X1  OAI21X1_30
timestamp 1560662619
transform -1 0 420 0 -1 505
box 0 0 32 100
use AOI21X1  AOI21X1_14
timestamp 1560662619
transform 1 0 420 0 -1 505
box 0 0 32 100
use FILL  FILL_4_0_0
timestamp 1560662619
transform 1 0 452 0 -1 505
box 0 0 8 100
use FILL  FILL_4_0_1
timestamp 1560662619
transform 1 0 460 0 -1 505
box 0 0 8 100
use OAI22X1  OAI22X1_4
timestamp 1560662619
transform 1 0 468 0 -1 505
box 0 0 40 100
use INVX2  INVX2_5
timestamp 1560662619
transform -1 0 524 0 -1 505
box 0 0 16 100
use NOR2X1  NOR2X1_33
timestamp 1560662619
transform 1 0 524 0 -1 505
box 0 0 24 100
use NOR2X1  NOR2X1_31
timestamp 1560662619
transform 1 0 548 0 -1 505
box 0 0 24 100
use AOI21X1  AOI21X1_16
timestamp 1560662619
transform 1 0 572 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_17
timestamp 1560662619
transform -1 0 636 0 -1 505
box 0 0 32 100
use INVX2  INVX2_4
timestamp 1560662619
transform 1 0 636 0 -1 505
box 0 0 16 100
use NOR2X1  NOR2X1_19
timestamp 1560662619
transform 1 0 652 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_34
timestamp 1560662619
transform 1 0 676 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_31
timestamp 1560662619
transform 1 0 700 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_1
timestamp 1560662619
transform 1 0 732 0 -1 505
box 0 0 24 100
use AND2X2  AND2X2_1
timestamp 1560662619
transform 1 0 756 0 -1 505
box 0 0 32 100
use INVX2  INVX2_3
timestamp 1560662619
transform 1 0 788 0 -1 505
box 0 0 16 100
use NAND2X1  NAND2X1_19
timestamp 1560662619
transform -1 0 828 0 -1 505
box 0 0 24 100
use OAI21X1  OAI21X1_29
timestamp 1560662619
transform 1 0 828 0 -1 505
box 0 0 32 100
use AOI21X1  AOI21X1_13
timestamp 1560662619
transform -1 0 892 0 -1 505
box 0 0 32 100
use OAI21X1  OAI21X1_9
timestamp 1560662619
transform -1 0 924 0 -1 505
box 0 0 32 100
use NOR2X1  NOR2X1_30
timestamp 1560662619
transform -1 0 948 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_38
timestamp 1560662619
transform 1 0 948 0 -1 505
box 0 0 24 100
use FILL  FILL_4_1_0
timestamp 1560662619
transform -1 0 980 0 -1 505
box 0 0 8 100
use FILL  FILL_4_1_1
timestamp 1560662619
transform -1 0 988 0 -1 505
box 0 0 8 100
use NOR2X1  NOR2X1_27
timestamp 1560662619
transform -1 0 1012 0 -1 505
box 0 0 24 100
use NAND3X1  NAND3X1_12
timestamp 1560662619
transform 1 0 1012 0 -1 505
box 0 0 32 100
use NOR2X1  NOR2X1_22
timestamp 1560662619
transform 1 0 1044 0 -1 505
box 0 0 24 100
use NAND3X1  NAND3X1_15
timestamp 1560662619
transform -1 0 1100 0 -1 505
box 0 0 32 100
use AOI21X1  AOI21X1_6
timestamp 1560662619
transform -1 0 1132 0 -1 505
box 0 0 32 100
use INVX1  INVX1_33
timestamp 1560662619
transform 1 0 1132 0 -1 505
box 0 0 16 100
use NAND2X1  NAND2X1_25
timestamp 1560662619
transform 1 0 1148 0 -1 505
box 0 0 24 100
use AOI21X1  AOI21X1_9
timestamp 1560662619
transform -1 0 1204 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_29
timestamp 1560662619
transform 1 0 1204 0 -1 505
box 0 0 24 100
use INVX2  INVX2_10
timestamp 1560662619
transform -1 0 1244 0 -1 505
box 0 0 16 100
use AOI21X1  AOI21X1_10
timestamp 1560662619
transform -1 0 1276 0 -1 505
box 0 0 32 100
use AOI21X1  AOI21X1_11
timestamp 1560662619
transform -1 0 1308 0 -1 505
box 0 0 32 100
use NOR2X1  NOR2X1_28
timestamp 1560662619
transform -1 0 1332 0 -1 505
box 0 0 24 100
use NOR2X1  NOR2X1_29
timestamp 1560662619
transform -1 0 1356 0 -1 505
box 0 0 24 100
use XNOR2X1  XNOR2X1_1
timestamp 1560662619
transform -1 0 1412 0 -1 505
box 0 0 56 100
use BUFX2  BUFX2_5
timestamp 1560662619
transform 1 0 1412 0 -1 505
box 0 0 24 100
use FILL  FILL_5_1
timestamp 1560662619
transform -1 0 1444 0 -1 505
box 0 0 8 100
use BUFX4  BUFX4_9
timestamp 1560662619
transform 1 0 4 0 1 305
box 0 0 32 100
use DFFSR  DFFSR_40
timestamp 1560662619
transform 1 0 36 0 1 305
box 0 0 176 100
use DFFSR  DFFSR_38
timestamp 1560662619
transform 1 0 212 0 1 305
box 0 0 176 100
use INVX2  INVX2_6
timestamp 1560662619
transform -1 0 404 0 1 305
box 0 0 16 100
use NAND2X1  NAND2X1_35
timestamp 1560662619
transform 1 0 404 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_1
timestamp 1560662619
transform 1 0 428 0 1 305
box 0 0 32 100
use FILL  FILL_3_0_0
timestamp 1560662619
transform 1 0 460 0 1 305
box 0 0 8 100
use FILL  FILL_3_0_1
timestamp 1560662619
transform 1 0 468 0 1 305
box 0 0 8 100
use AOI21X1  AOI21X1_20
timestamp 1560662619
transform 1 0 476 0 1 305
box 0 0 32 100
use INVX1  INVX1_37
timestamp 1560662619
transform 1 0 508 0 1 305
box 0 0 16 100
use OAI21X1  OAI21X1_32
timestamp 1560662619
transform 1 0 524 0 1 305
box 0 0 32 100
use NAND3X1  NAND3X1_19
timestamp 1560662619
transform -1 0 588 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_32
timestamp 1560662619
transform 1 0 588 0 1 305
box 0 0 24 100
use AOI22X1  AOI22X1_3
timestamp 1560662619
transform -1 0 652 0 1 305
box 0 0 40 100
use NAND2X1  NAND2X1_21
timestamp 1560662619
transform -1 0 676 0 1 305
box 0 0 24 100
use AOI21X1  AOI21X1_18
timestamp 1560662619
transform -1 0 708 0 1 305
box 0 0 32 100
use INVX1  INVX1_36
timestamp 1560662619
transform 1 0 708 0 1 305
box 0 0 16 100
use AOI21X1  AOI21X1_17
timestamp 1560662619
transform -1 0 756 0 1 305
box 0 0 32 100
use NAND3X1  NAND3X1_18
timestamp 1560662619
transform -1 0 788 0 1 305
box 0 0 32 100
use AOI22X1  AOI22X1_2
timestamp 1560662619
transform -1 0 828 0 1 305
box 0 0 40 100
use AOI21X1  AOI21X1_15
timestamp 1560662619
transform -1 0 860 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_20
timestamp 1560662619
transform 1 0 860 0 1 305
box 0 0 24 100
use OAI21X1  OAI21X1_11
timestamp 1560662619
transform 1 0 884 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_31
timestamp 1560662619
transform -1 0 940 0 1 305
box 0 0 24 100
use INVX2  INVX2_2
timestamp 1560662619
transform -1 0 956 0 1 305
box 0 0 16 100
use FILL  FILL_3_1_0
timestamp 1560662619
transform 1 0 956 0 1 305
box 0 0 8 100
use FILL  FILL_3_1_1
timestamp 1560662619
transform 1 0 964 0 1 305
box 0 0 8 100
use BUFX4  BUFX4_7
timestamp 1560662619
transform 1 0 972 0 1 305
box 0 0 32 100
use NAND3X1  NAND3X1_16
timestamp 1560662619
transform 1 0 1004 0 1 305
box 0 0 32 100
use OAI22X1  OAI22X1_3
timestamp 1560662619
transform -1 0 1076 0 1 305
box 0 0 40 100
use INVX8  INVX8_2
timestamp 1560662619
transform 1 0 1076 0 1 305
box 0 0 40 100
use INVX4  INVX4_2
timestamp 1560662619
transform 1 0 1116 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_27
timestamp 1560662619
transform 1 0 1140 0 1 305
box 0 0 24 100
use OAI21X1  OAI21X1_26
timestamp 1560662619
transform -1 0 1196 0 1 305
box 0 0 32 100
use AOI21X1  AOI21X1_7
timestamp 1560662619
transform 1 0 1196 0 1 305
box 0 0 32 100
use DFFSR  DFFSR_12
timestamp 1560662619
transform -1 0 1404 0 1 305
box 0 0 176 100
use BUFX2  BUFX2_4
timestamp 1560662619
transform 1 0 1404 0 1 305
box 0 0 24 100
use FILL  FILL_4_1
timestamp 1560662619
transform 1 0 1428 0 1 305
box 0 0 8 100
use FILL  FILL_4_2
timestamp 1560662619
transform 1 0 1436 0 1 305
box 0 0 8 100
use DFFSR  DFFSR_35
timestamp 1560662619
transform 1 0 4 0 -1 305
box 0 0 176 100
use DFFSR  DFFSR_41
timestamp 1560662619
transform 1 0 180 0 -1 305
box 0 0 176 100
use INVX2  INVX2_7
timestamp 1560662619
transform 1 0 356 0 -1 305
box 0 0 16 100
use NOR2X1  NOR2X1_36
timestamp 1560662619
transform -1 0 396 0 -1 305
box 0 0 24 100
use OAI22X1  OAI22X1_5
timestamp 1560662619
transform 1 0 396 0 -1 305
box 0 0 40 100
use NOR2X1  NOR2X1_34
timestamp 1560662619
transform -1 0 460 0 -1 305
box 0 0 24 100
use FILL  FILL_2_0_0
timestamp 1560662619
transform 1 0 460 0 -1 305
box 0 0 8 100
use FILL  FILL_2_0_1
timestamp 1560662619
transform 1 0 468 0 -1 305
box 0 0 8 100
use AOI21X1  AOI21X1_19
timestamp 1560662619
transform 1 0 476 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_20
timestamp 1560662619
transform 1 0 508 0 -1 305
box 0 0 24 100
use INVX1  INVX1_24
timestamp 1560662619
transform 1 0 532 0 -1 305
box 0 0 16 100
use OAI21X1  OAI21X1_14
timestamp 1560662619
transform 1 0 548 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_35
timestamp 1560662619
transform -1 0 604 0 -1 305
box 0 0 24 100
use NOR2X1  NOR2X1_1
timestamp 1560662619
transform 1 0 604 0 -1 305
box 0 0 24 100
use OAI21X1  OAI21X1_13
timestamp 1560662619
transform 1 0 628 0 -1 305
box 0 0 32 100
use BUFX4  BUFX4_14
timestamp 1560662619
transform 1 0 660 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_8
timestamp 1560662619
transform 1 0 692 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_33
timestamp 1560662619
transform 1 0 724 0 -1 305
box 0 0 24 100
use BUFX4  BUFX4_1
timestamp 1560662619
transform 1 0 748 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_24
timestamp 1560662619
transform 1 0 780 0 -1 305
box 0 0 24 100
use NAND2X1  NAND2X1_30
timestamp 1560662619
transform 1 0 804 0 -1 305
box 0 0 24 100
use AOI21X1  AOI21X1_12
timestamp 1560662619
transform -1 0 860 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_7
timestamp 1560662619
transform -1 0 892 0 -1 305
box 0 0 32 100
use NAND3X1  NAND3X1_13
timestamp 1560662619
transform -1 0 924 0 -1 305
box 0 0 32 100
use INVX1  INVX1_34
timestamp 1560662619
transform 1 0 924 0 -1 305
box 0 0 16 100
use NAND3X1  NAND3X1_14
timestamp 1560662619
transform 1 0 940 0 -1 305
box 0 0 32 100
use FILL  FILL_2_1_0
timestamp 1560662619
transform 1 0 972 0 -1 305
box 0 0 8 100
use FILL  FILL_2_1_1
timestamp 1560662619
transform 1 0 980 0 -1 305
box 0 0 8 100
use NAND2X1  NAND2X1_16
timestamp 1560662619
transform 1 0 988 0 -1 305
box 0 0 24 100
use DFFSR  DFFSR_34
timestamp 1560662619
transform -1 0 1188 0 -1 305
box 0 0 176 100
use DFFSR  DFFSR_13
timestamp 1560662619
transform -1 0 1364 0 -1 305
box 0 0 176 100
use CLKBUF1  CLKBUF1_6
timestamp 1560662619
transform -1 0 1436 0 -1 305
box 0 0 72 100
use FILL  FILL_3_1
timestamp 1560662619
transform -1 0 1444 0 -1 305
box 0 0 8 100
use CLKBUF1  CLKBUF1_5
timestamp 1560662619
transform 1 0 4 0 1 105
box 0 0 72 100
use DFFSR  DFFSR_42
timestamp 1560662619
transform 1 0 76 0 1 105
box 0 0 176 100
use NOR3X1  NOR3X1_8
timestamp 1560662619
transform -1 0 316 0 1 105
box 0 0 64 100
use NAND2X1  NAND2X1_36
timestamp 1560662619
transform 1 0 316 0 1 105
box 0 0 24 100
use AND2X2  AND2X2_5
timestamp 1560662619
transform 1 0 340 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_33
timestamp 1560662619
transform 1 0 372 0 1 105
box 0 0 32 100
use INVX2  INVX2_8
timestamp 1560662619
transform -1 0 420 0 1 105
box 0 0 16 100
use AOI21X1  AOI21X1_21
timestamp 1560662619
transform -1 0 452 0 1 105
box 0 0 32 100
use FILL  FILL_1_0_0
timestamp 1560662619
transform -1 0 460 0 1 105
box 0 0 8 100
use FILL  FILL_1_0_1
timestamp 1560662619
transform -1 0 468 0 1 105
box 0 0 8 100
use AOI22X1  AOI22X1_4
timestamp 1560662619
transform -1 0 508 0 1 105
box 0 0 40 100
use NAND2X1  NAND2X1_23
timestamp 1560662619
transform -1 0 532 0 1 105
box 0 0 24 100
use AOI21X1  AOI21X1_22
timestamp 1560662619
transform 1 0 532 0 1 105
box 0 0 32 100
use NAND2X1  NAND2X1_22
timestamp 1560662619
transform -1 0 588 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_15
timestamp 1560662619
transform -1 0 620 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_2
timestamp 1560662619
transform 1 0 620 0 1 105
box 0 0 24 100
use BUFX4  BUFX4_11
timestamp 1560662619
transform 1 0 644 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_13
timestamp 1560662619
transform 1 0 676 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_2
timestamp 1560662619
transform 1 0 708 0 1 105
box 0 0 32 100
use BUFX4  BUFX4_3
timestamp 1560662619
transform 1 0 740 0 1 105
box 0 0 32 100
use INVX8  INVX8_3
timestamp 1560662619
transform -1 0 812 0 1 105
box 0 0 40 100
use NOR2X1  NOR2X1_17
timestamp 1560662619
transform 1 0 812 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_18
timestamp 1560662619
transform 1 0 836 0 1 105
box 0 0 24 100
use NOR2X1  NOR2X1_21
timestamp 1560662619
transform 1 0 860 0 1 105
box 0 0 24 100
use AOI21X1  AOI21X1_5
timestamp 1560662619
transform -1 0 916 0 1 105
box 0 0 32 100
use AOI21X1  AOI21X1_8
timestamp 1560662619
transform -1 0 948 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_22
timestamp 1560662619
transform -1 0 980 0 1 105
box 0 0 32 100
use FILL  FILL_1_1_0
timestamp 1560662619
transform -1 0 988 0 1 105
box 0 0 8 100
use FILL  FILL_1_1_1
timestamp 1560662619
transform -1 0 996 0 1 105
box 0 0 8 100
use OAI21X1  OAI21X1_21
timestamp 1560662619
transform -1 0 1028 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_16
timestamp 1560662619
transform -1 0 1052 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_18
timestamp 1560662619
transform -1 0 1084 0 1 105
box 0 0 32 100
use NOR2X1  NOR2X1_23
timestamp 1560662619
transform -1 0 1108 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_19
timestamp 1560662619
transform 1 0 1108 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_3
timestamp 1560662619
transform 1 0 1140 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_20
timestamp 1560662619
transform 1 0 1172 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_17
timestamp 1560662619
transform 1 0 1204 0 1 105
box 0 0 32 100
use INVX1  INVX1_11
timestamp 1560662619
transform -1 0 1252 0 1 105
box 0 0 16 100
use DFFSR  DFFSR_14
timestamp 1560662619
transform -1 0 1428 0 1 105
box 0 0 176 100
use FILL  FILL_2_1
timestamp 1560662619
transform 1 0 1428 0 1 105
box 0 0 8 100
use FILL  FILL_2_2
timestamp 1560662619
transform 1 0 1436 0 1 105
box 0 0 8 100
use BUFX2  BUFX2_19
timestamp 1560662619
transform 1 0 4 0 -1 105
box 0 0 24 100
use CLKBUF1  CLKBUF1_2
timestamp 1560662619
transform 1 0 28 0 -1 105
box 0 0 72 100
use DFFSR  DFFSR_43
timestamp 1560662619
transform 1 0 100 0 -1 105
box 0 0 176 100
use NOR2X1  NOR2X1_38
timestamp 1560662619
transform 1 0 276 0 -1 105
box 0 0 24 100
use AOI21X1  AOI21X1_25
timestamp 1560662619
transform -1 0 332 0 -1 105
box 0 0 32 100
use NOR3X1  NOR3X1_9
timestamp 1560662619
transform 1 0 332 0 -1 105
box 0 0 64 100
use OAI21X1  OAI21X1_34
timestamp 1560662619
transform -1 0 428 0 -1 105
box 0 0 32 100
use INVX1  INVX1_25
timestamp 1560662619
transform 1 0 428 0 -1 105
box 0 0 16 100
use FILL  FILL_0_0_0
timestamp 1560662619
transform 1 0 444 0 -1 105
box 0 0 8 100
use FILL  FILL_0_0_1
timestamp 1560662619
transform 1 0 452 0 -1 105
box 0 0 8 100
use AOI21X1  AOI21X1_23
timestamp 1560662619
transform 1 0 460 0 -1 105
box 0 0 32 100
use AOI21X1  AOI21X1_24
timestamp 1560662619
transform -1 0 524 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_16
timestamp 1560662619
transform 1 0 524 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_6
timestamp 1560662619
transform -1 0 588 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_37
timestamp 1560662619
transform -1 0 612 0 -1 105
box 0 0 24 100
use NOR2X1  NOR2X1_37
timestamp 1560662619
transform 1 0 612 0 -1 105
box 0 0 24 100
use BUFX4  BUFX4_12
timestamp 1560662619
transform -1 0 668 0 -1 105
box 0 0 32 100
use BUFX4  BUFX4_4
timestamp 1560662619
transform -1 0 700 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_17
timestamp 1560662619
transform 1 0 700 0 -1 105
box 0 0 24 100
use DFFSR  DFFSR_33
timestamp 1560662619
transform -1 0 900 0 -1 105
box 0 0 176 100
use NOR2X1  NOR2X1_24
timestamp 1560662619
transform -1 0 924 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_26
timestamp 1560662619
transform -1 0 948 0 -1 105
box 0 0 24 100
use OAI21X1  OAI21X1_23
timestamp 1560662619
transform 1 0 948 0 -1 105
box 0 0 32 100
use FILL  FILL_0_1_0
timestamp 1560662619
transform -1 0 988 0 -1 105
box 0 0 8 100
use FILL  FILL_0_1_1
timestamp 1560662619
transform -1 0 996 0 -1 105
box 0 0 8 100
use AND2X2  AND2X2_4
timestamp 1560662619
transform -1 0 1028 0 -1 105
box 0 0 32 100
use INVX1  INVX1_10
timestamp 1560662619
transform -1 0 1044 0 -1 105
box 0 0 16 100
use INVX1  INVX1_35
timestamp 1560662619
transform 1 0 1044 0 -1 105
box 0 0 16 100
use OAI21X1  OAI21X1_24
timestamp 1560662619
transform 1 0 1060 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_25
timestamp 1560662619
transform -1 0 1124 0 -1 105
box 0 0 32 100
use NOR2X1  NOR2X1_25
timestamp 1560662619
transform -1 0 1148 0 -1 105
box 0 0 24 100
use DFFSR  DFFSR_15
timestamp 1560662619
transform -1 0 1324 0 -1 105
box 0 0 176 100
use INVX1  INVX1_15
timestamp 1560662619
transform -1 0 1340 0 -1 105
box 0 0 16 100
use BUFX2  BUFX2_3
timestamp 1560662619
transform 1 0 1340 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_16
timestamp 1560662619
transform -1 0 1388 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_10
timestamp 1560662619
transform 1 0 1388 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_14
timestamp 1560662619
transform -1 0 1436 0 -1 105
box 0 0 24 100
use FILL  FILL_1_1
timestamp 1560662619
transform -1 0 1444 0 -1 105
box 0 0 8 100
use PADINC  PADINC_1
timestamp 1560662619
transform 0 1 1666 -1 0 1548
box 0 0 900 3000
use PADINC  PADINC_3
timestamp 1560662619
transform 0 -1 -98 1 0 -240
box 0 0 900 3000
use PADFC  PADFC_3
timestamp 1560662619
transform 1 0 -3098 0 -1 -228
box 0 0 3000 3000
use PADINC  PADINC_0
timestamp 1560662619
transform -1 0 790 0 -1 -228
box 0 0 900 3000
use PADOUT  PADOUT_0
timestamp 1560662619
transform 0 1 1666 -1 0 660
box 0 0 900 3000
use PADGND  PADGND_1
timestamp 1560662619
transform -1 0 1678 0 -1 -228
box 0 0 900 3000
use PADFC  PADFC_2
timestamp 1560662619
transform -1 0 4666 0 -1 -228
box 0 0 3000 3000
<< labels >>
rlabel metal6 440 -30 456 -22 8 vdd
port 0 nsew
rlabel metal6 960 -30 976 -22 8 gnd
port 1 nsew
rlabel metal3 -26 1288 -22 1292 4 RST
port 2 nsew
rlabel metal3 -26 138 -22 142 4 SCK
port 3 nsew
rlabel metal3 -26 558 -22 562 4 SDI
port 4 nsew
rlabel metal3 -26 1248 -22 1252 4 CSB
port 5 nsew
rlabel metal3 1470 1318 1474 1322 6 trap
port 6 nsew
rlabel metal2 1310 -22 1314 -18 8 mask_rev_in[0]
port 7 nsew
rlabel metal2 1406 -22 1410 -18 8 mask_rev_in[1]
port 8 nsew
rlabel metal2 1422 -22 1426 -18 8 mask_rev_in[2]
port 9 nsew
rlabel metal2 1438 -22 1442 -18 8 mask_rev_in[3]
port 10 nsew
rlabel metal3 -26 1308 -22 1312 4 SDO
port 11 nsew
rlabel metal3 -26 1148 -22 1152 4 sdo_enb
port 12 nsew
rlabel metal3 -26 1268 -22 1272 4 xtal_ena
port 13 nsew
rlabel metal2 1014 1328 1018 1332 6 reg_ena
port 14 nsew
rlabel metal2 1302 1328 1306 1332 6 pll_vco_ena
port 15 nsew
rlabel metal2 998 1328 1002 1332 6 pll_cp_ena
port 16 nsew
rlabel metal2 14 -22 18 -18 8 pll_bias_ena
port 17 nsew
rlabel metal2 934 1328 938 1332 6 pll_trim[0]
port 18 nsew
rlabel metal2 486 1328 490 1332 6 pll_trim[1]
port 19 nsew
rlabel metal2 270 1328 274 1332 6 pll_trim[2]
port 20 nsew
rlabel metal2 62 1328 66 1332 6 pll_trim[3]
port 21 nsew
rlabel metal3 1470 1258 1474 1262 6 pll_bypass
port 22 nsew
rlabel metal3 1470 1278 1474 1282 6 irq
port 23 nsew
rlabel metal3 1470 1298 1474 1302 6 reset
port 24 nsew
rlabel metal3 1470 1018 1474 1022 6 mfgr_id[0]
port 25 nsew
rlabel metal3 1470 1038 1474 1042 6 mfgr_id[1]
port 26 nsew
rlabel metal3 1470 1058 1474 1062 6 mfgr_id[2]
port 27 nsew
rlabel metal3 1470 1078 1474 1082 6 mfgr_id[3]
port 28 nsew
rlabel metal3 1470 1098 1474 1102 6 mfgr_id[4]
port 29 nsew
rlabel metal3 1470 1118 1474 1122 6 mfgr_id[5]
port 30 nsew
rlabel metal3 1470 1138 1474 1142 6 mfgr_id[6]
port 31 nsew
rlabel metal3 1470 1158 1474 1162 6 mfgr_id[7]
port 32 nsew
rlabel metal3 1470 1178 1474 1182 6 mfgr_id[8]
port 33 nsew
rlabel metal3 1470 1198 1474 1202 6 mfgr_id[9]
port 34 nsew
rlabel metal3 1470 1218 1474 1222 6 mfgr_id[10]
port 35 nsew
rlabel metal3 1470 1238 1474 1242 6 mfgr_id[11]
port 36 nsew
rlabel metal2 1318 1328 1322 1332 6 prod_id[0]
port 37 nsew
rlabel metal2 1334 1328 1338 1332 6 prod_id[1]
port 38 nsew
rlabel metal2 1350 1328 1354 1332 6 prod_id[2]
port 39 nsew
rlabel metal2 1366 1328 1370 1332 6 prod_id[3]
port 40 nsew
rlabel metal2 1382 1328 1386 1332 6 prod_id[4]
port 41 nsew
rlabel metal2 1398 1328 1402 1332 6 prod_id[5]
port 42 nsew
rlabel metal2 1414 1328 1418 1332 6 prod_id[6]
port 43 nsew
rlabel metal2 1430 1328 1434 1332 6 prod_id[7]
port 44 nsew
rlabel metal3 1470 48 1474 52 6 mask_rev[0]
port 45 nsew
rlabel metal3 1470 348 1474 352 6 mask_rev[1]
port 46 nsew
rlabel metal3 1470 448 1474 452 6 mask_rev[2]
port 47 nsew
rlabel metal3 1470 648 1474 652 6 mask_rev[3]
port 48 nsew
<< end >>
